module attack_FSM (
    input logic btn_atk,
    input logic btn_up,
    input logic btn_down,
    input logic btn_right,
    input logic btn_left,
    input logic hit_stun_active,
    output logic attack_active,
    output logic anim_ID,
);
//always_comb begin
//if (hit_stun_active) 
//end

endmodule