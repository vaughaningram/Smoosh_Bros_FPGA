module ROM_Screen (
    input logic clk,
    input logic [16:0] addr,
    output logic [5:0] data
    // logic timer = counter[25]; // timer for changing addresses. Depends on what
    //                         // speed you need. 
);


logic [5:0] data_comb;
// // HSOSC component -> On chip oscillator
//     SB_HFOSC #(
//         .CLKHF_DIV("0b00")
//     ) osc (
//         .CLKHFPU(1'b1), // Power up
//         .CLKHFEN(1'b1), // Enable
//         .CLKHF(clk)     // Clock output
//         // (TRIM pins omitted intentionally)
//     );

always_ff @(posedge clk) begin
    data <= data_comb; // takes data from ROM on clock tick to data
end

// always_ff @(posedge timer) begin
//     addr <= addr + 1; // increment address
// end

// writing always_comb in this way tells System Verilog it is ROM
always_comb begin
    case(addr)
  17'b00000000000000000 : data_comb = 6'b000101;
 17'b00000000000000001 : data_comb = 6'b000101;
 17'b00000000000000010 : data_comb = 6'b000101;
 17'b00000000000000011 : data_comb = 6'b000101;
 17'b00000000000000100 : data_comb = 6'b000101;
 17'b00000000000000101 : data_comb = 6'b000101;
 17'b00000000000000110 : data_comb = 6'b000101;
 17'b00000000000000111 : data_comb = 6'b000101;
 17'b00000000000001000 : data_comb = 6'b000101;
 17'b00000000000001001 : data_comb = 6'b000101;
 17'b00000000000001010 : data_comb = 6'b000101;
 17'b00000000000001011 : data_comb = 6'b000101;
 17'b00000000000001100 : data_comb = 6'b000101;
 17'b00000000000001101 : data_comb = 6'b000101;
 17'b00000000000001110 : data_comb = 6'b000101;
 17'b00000000000001111 : data_comb = 6'b000101;
 17'b00000000000010000 : data_comb = 6'b000101;
 17'b00000000000010001 : data_comb = 6'b000101;
 17'b00000000000010010 : data_comb = 6'b000101;
 17'b00000000000010011 : data_comb = 6'b000101;
 17'b00000000000010100 : data_comb = 6'b000101;
 17'b00000000000010101 : data_comb = 6'b000101;
 17'b00000000000010110 : data_comb = 6'b000101;
 17'b00000000000010111 : data_comb = 6'b000101;
 17'b00000000000011000 : data_comb = 6'b000101;
 17'b00000000000011001 : data_comb = 6'b000101;
 17'b00000000000011010 : data_comb = 6'b000101;
 17'b00000000000011011 : data_comb = 6'b000101;
 17'b00000000000011100 : data_comb = 6'b000101;
 17'b00000000000011101 : data_comb = 6'b000101;
 17'b00000000000011110 : data_comb = 6'b000101;
 17'b00000000000011111 : data_comb = 6'b000101;
 17'b00000000000100000 : data_comb = 6'b000101;
 17'b00000000000100001 : data_comb = 6'b000101;
 17'b00000000000100010 : data_comb = 6'b000101;
 17'b00000000000100011 : data_comb = 6'b000101;
 17'b00000000000100100 : data_comb = 6'b000101;
 17'b00000000000100101 : data_comb = 6'b000101;
 17'b00000000000100110 : data_comb = 6'b000101;
 17'b00000000000100111 : data_comb = 6'b000101;
 17'b00000000000101000 : data_comb = 6'b000101;
 17'b00000000000101001 : data_comb = 6'b000101;
 17'b00000000000101010 : data_comb = 6'b000101;
 17'b00000000000101011 : data_comb = 6'b000101;
 17'b00000000000101100 : data_comb = 6'b000101;
 17'b00000000000101101 : data_comb = 6'b000101;
 17'b00000000000101110 : data_comb = 6'b000101;
 17'b00000000000101111 : data_comb = 6'b000101;
 17'b00000000000110000 : data_comb = 6'b000101;
 17'b00000000000110001 : data_comb = 6'b000101;
 17'b00000000000110010 : data_comb = 6'b000101;
 17'b00000000000110011 : data_comb = 6'b000101;
 17'b00000000000110100 : data_comb = 6'b000101;
 17'b00000000000110101 : data_comb = 6'b000101;
 17'b00000000000110110 : data_comb = 6'b000101;
 17'b00000000000110111 : data_comb = 6'b000101;
 17'b00000000000111000 : data_comb = 6'b000101;
 17'b00000000000111001 : data_comb = 6'b000101;
 17'b00000000000111010 : data_comb = 6'b000101;
 17'b00000000000111011 : data_comb = 6'b000101;
 17'b00000000000111100 : data_comb = 6'b000101;
 17'b00000000000111101 : data_comb = 6'b000101;
 17'b00000000000111110 : data_comb = 6'b000101;
 17'b00000000000111111 : data_comb = 6'b000101;
 17'b00000000001000000 : data_comb = 6'b000101;
 17'b00000000001000001 : data_comb = 6'b000101;
 17'b00000000001000010 : data_comb = 6'b000101;
 17'b00000000001000011 : data_comb = 6'b000101;
 17'b00000000001000100 : data_comb = 6'b000101;
 17'b00000000001000101 : data_comb = 6'b000101;
 17'b00000000001000110 : data_comb = 6'b000101;
 17'b00000000001000111 : data_comb = 6'b000101;
 17'b00000000001001000 : data_comb = 6'b000101;
 17'b00000000001001001 : data_comb = 6'b000101;
 17'b00000000001001010 : data_comb = 6'b000101;
 17'b00000000001001011 : data_comb = 6'b000101;
 17'b00000000001001100 : data_comb = 6'b000101;
 17'b00000000001001101 : data_comb = 6'b000101;
 17'b00000000001001110 : data_comb = 6'b000101;
 17'b00000000001001111 : data_comb = 6'b000101;
 17'b00000000001010000 : data_comb = 6'b000101;
 17'b00000000001010001 : data_comb = 6'b000101;
 17'b00000000001010010 : data_comb = 6'b000101;
 17'b00000000001010011 : data_comb = 6'b000101;
 17'b00000000001010100 : data_comb = 6'b000101;
 17'b00000000001010101 : data_comb = 6'b000101;
 17'b00000000001010110 : data_comb = 6'b000101;
 17'b00000000001010111 : data_comb = 6'b000101;
 17'b00000000001011000 : data_comb = 6'b000101;
 17'b00000000001011001 : data_comb = 6'b000101;
 17'b00000000001011010 : data_comb = 6'b000101;
 17'b00000000001011011 : data_comb = 6'b000101;
 17'b00000000001011100 : data_comb = 6'b000101;
 17'b00000000001011101 : data_comb = 6'b000101;
 17'b00000000001011110 : data_comb = 6'b000101;
 17'b00000000001011111 : data_comb = 6'b000101;
 17'b00000000001100000 : data_comb = 6'b000101;
 17'b00000000001100001 : data_comb = 6'b000101;
 17'b00000000001100010 : data_comb = 6'b000101;
 17'b00000000001100011 : data_comb = 6'b000101;
 17'b00000000001100100 : data_comb = 6'b000101;
 17'b00000000001100101 : data_comb = 6'b000101;
 17'b00000000001100110 : data_comb = 6'b000101;
 17'b00000000001100111 : data_comb = 6'b000101;
 17'b00000000001101000 : data_comb = 6'b000101;
 17'b00000000001101001 : data_comb = 6'b000101;
 17'b00000000001101010 : data_comb = 6'b000101;
 17'b00000000001101011 : data_comb = 6'b000101;
 17'b00000000001101100 : data_comb = 6'b000101;
 17'b00000000001101101 : data_comb = 6'b000101;
 17'b00000000001101110 : data_comb = 6'b000101;
 17'b00000000001101111 : data_comb = 6'b000101;
 17'b00000000001110000 : data_comb = 6'b000101;
 17'b00000000001110001 : data_comb = 6'b000101;
 17'b00000000001110010 : data_comb = 6'b000101;
 17'b00000000001110011 : data_comb = 6'b000101;
 17'b00000000001110100 : data_comb = 6'b000101;
 17'b00000000001110101 : data_comb = 6'b000101;
 17'b00000000001110110 : data_comb = 6'b000101;
 17'b00000000001110111 : data_comb = 6'b000101;
 17'b00000000001111000 : data_comb = 6'b000101;
 17'b00000000001111001 : data_comb = 6'b000101;
 17'b00000000001111010 : data_comb = 6'b000101;
 17'b00000000001111011 : data_comb = 6'b000101;
 17'b00000000001111100 : data_comb = 6'b000101;
 17'b00000000001111101 : data_comb = 6'b000101;
 17'b00000000001111110 : data_comb = 6'b000101;
 17'b00000000001111111 : data_comb = 6'b000101;
 17'b00000000010000000 : data_comb = 6'b000101;
 17'b00000000010000001 : data_comb = 6'b000101;
 17'b00000000010000010 : data_comb = 6'b000101;
 17'b00000000010000011 : data_comb = 6'b000101;
 17'b00000000010000100 : data_comb = 6'b000101;
 17'b00000000010000101 : data_comb = 6'b000101;
 17'b00000000010000110 : data_comb = 6'b000101;
 17'b00000000010000111 : data_comb = 6'b000101;
 17'b00000000010001000 : data_comb = 6'b000101;
 17'b00000000010001001 : data_comb = 6'b000101;
 17'b00000000010001010 : data_comb = 6'b000101;
 17'b00000000010001011 : data_comb = 6'b000101;
 17'b00000000010001100 : data_comb = 6'b000101;
 17'b00000000010001101 : data_comb = 6'b000101;
 17'b00000000010001110 : data_comb = 6'b000101;
 17'b00000000010001111 : data_comb = 6'b000101;
 17'b00000000010010000 : data_comb = 6'b000101;
 17'b00000000010010001 : data_comb = 6'b000101;
 17'b00000000010010010 : data_comb = 6'b000101;
 17'b00000000010010011 : data_comb = 6'b000101;
 17'b00000000010010100 : data_comb = 6'b000101;
 17'b00000000010010101 : data_comb = 6'b000101;
 17'b00000000010010110 : data_comb = 6'b000101;
 17'b00000000010010111 : data_comb = 6'b000101;
 17'b00000000010011000 : data_comb = 6'b000101;
 17'b00000000010011001 : data_comb = 6'b000101;
 17'b00000000010011010 : data_comb = 6'b000101;
 17'b00000000010011011 : data_comb = 6'b000101;
 17'b00000000010011100 : data_comb = 6'b000101;
 17'b00000000010011101 : data_comb = 6'b000101;
 17'b00000000010011110 : data_comb = 6'b000101;
 17'b00000000010011111 : data_comb = 6'b000101;
 17'b00000000010100000 : data_comb = 6'b000101;
 17'b00000000010100001 : data_comb = 6'b000101;
 17'b00000000010100010 : data_comb = 6'b000101;
 17'b00000000010100011 : data_comb = 6'b000101;
 17'b00000000010100100 : data_comb = 6'b000101;
 17'b00000000010100101 : data_comb = 6'b000101;
 17'b00000000010100110 : data_comb = 6'b000101;
 17'b00000000010100111 : data_comb = 6'b000101;
 17'b00000000010101000 : data_comb = 6'b000101;
 17'b00000000010101001 : data_comb = 6'b000101;
 17'b00000000010101010 : data_comb = 6'b000101;
 17'b00000000010101011 : data_comb = 6'b000101;
 17'b00000000010101100 : data_comb = 6'b000101;
 17'b00000000010101101 : data_comb = 6'b000101;
 17'b00000000010101110 : data_comb = 6'b000101;
 17'b00000000010101111 : data_comb = 6'b000101;
 17'b00000000010110000 : data_comb = 6'b000101;
 17'b00000000010110001 : data_comb = 6'b000101;
 17'b00000000010110010 : data_comb = 6'b000101;
 17'b00000000010110011 : data_comb = 6'b000101;
 17'b00000000010110100 : data_comb = 6'b000101;
 17'b00000000010110101 : data_comb = 6'b000101;
 17'b00000000010110110 : data_comb = 6'b000101;
 17'b00000000010110111 : data_comb = 6'b000101;
 17'b00000000010111000 : data_comb = 6'b000101;
 17'b00000000010111001 : data_comb = 6'b000101;
 17'b00000000010111010 : data_comb = 6'b000101;
 17'b00000000010111011 : data_comb = 6'b000101;
 17'b00000000010111100 : data_comb = 6'b000101;
 17'b00000000010111101 : data_comb = 6'b000101;
 17'b00000000010111110 : data_comb = 6'b000101;
 17'b00000000010111111 : data_comb = 6'b000101;
 17'b00000000011000000 : data_comb = 6'b000101;
 17'b00000000011000001 : data_comb = 6'b000101;
 17'b00000000011000010 : data_comb = 6'b000101;
 17'b00000000011000011 : data_comb = 6'b000101;
 17'b00000000011000100 : data_comb = 6'b000101;
 17'b00000000011000101 : data_comb = 6'b000101;
 17'b00000000011000110 : data_comb = 6'b000101;
 17'b00000000011000111 : data_comb = 6'b000101;
 17'b00000000011001000 : data_comb = 6'b000101;
 17'b00000000011001001 : data_comb = 6'b000101;
 17'b00000000011001010 : data_comb = 6'b000101;
 17'b00000000011001011 : data_comb = 6'b000101;
 17'b00000000011001100 : data_comb = 6'b000101;
 17'b00000000011001101 : data_comb = 6'b000101;
 17'b00000000011001110 : data_comb = 6'b000101;
 17'b00000000011001111 : data_comb = 6'b000101;
 17'b00000000011010000 : data_comb = 6'b000101;
 17'b00000000011010001 : data_comb = 6'b000101;
 17'b00000000011010010 : data_comb = 6'b000101;
 17'b00000000011010011 : data_comb = 6'b000101;
 17'b00000000011010100 : data_comb = 6'b000101;
 17'b00000000011010101 : data_comb = 6'b000101;
 17'b00000000011010110 : data_comb = 6'b000101;
 17'b00000000011010111 : data_comb = 6'b000101;
 17'b00000000011011000 : data_comb = 6'b000101;
 17'b00000000011011001 : data_comb = 6'b000101;
 17'b00000000011011010 : data_comb = 6'b000101;
 17'b00000000011011011 : data_comb = 6'b000101;
 17'b00000000011011100 : data_comb = 6'b000101;
 17'b00000000011011101 : data_comb = 6'b000101;
 17'b00000000011011110 : data_comb = 6'b000101;
 17'b00000000011011111 : data_comb = 6'b000101;
 17'b00000000011100000 : data_comb = 6'b000101;
 17'b00000000011100001 : data_comb = 6'b000101;
 17'b00000000011100010 : data_comb = 6'b000101;
 17'b00000000011100011 : data_comb = 6'b000101;
 17'b00000000011100100 : data_comb = 6'b000101;
 17'b00000000011100101 : data_comb = 6'b000101;
 17'b00000000011100110 : data_comb = 6'b000101;
 17'b00000000011100111 : data_comb = 6'b000101;
 17'b00000000011101000 : data_comb = 6'b000101;
 17'b00000000011101001 : data_comb = 6'b000101;
 17'b00000000011101010 : data_comb = 6'b000101;
 17'b00000000011101011 : data_comb = 6'b000101;
 17'b00000000011101100 : data_comb = 6'b000101;
 17'b00000000011101101 : data_comb = 6'b000101;
 17'b00000000011101110 : data_comb = 6'b000101;
 17'b00000000011101111 : data_comb = 6'b000101;
 17'b00000000011110000 : data_comb = 6'b000101;
 17'b00000000011110001 : data_comb = 6'b000101;
 17'b00000000011110010 : data_comb = 6'b000101;
 17'b00000000011110011 : data_comb = 6'b000101;
 17'b00000000011110100 : data_comb = 6'b000101;
 17'b00000000011110101 : data_comb = 6'b000101;
 17'b00000000011110110 : data_comb = 6'b000101;
 17'b00000000011110111 : data_comb = 6'b000101;
 17'b00000000011111000 : data_comb = 6'b000101;
 17'b00000000011111001 : data_comb = 6'b000101;
 17'b00000000011111010 : data_comb = 6'b000101;
 17'b00000000011111011 : data_comb = 6'b000101;
 17'b00000000011111100 : data_comb = 6'b010101;
 17'b00000000011111101 : data_comb = 6'b101000;
 17'b00000000011111110 : data_comb = 6'b101000;
 17'b00000000011111111 : data_comb = 6'b000101;
 17'b00000000100000000 : data_comb = 6'b000101;
 17'b00000000100000001 : data_comb = 6'b000101;
 17'b00000000100000010 : data_comb = 6'b000101;
 17'b00000000100000011 : data_comb = 6'b000101;
 17'b00000000100000100 : data_comb = 6'b000101;
 17'b00000000100000101 : data_comb = 6'b000101;
 17'b00000000100000110 : data_comb = 6'b000101;
 17'b00000000100000111 : data_comb = 6'b000101;
 17'b00000000100001000 : data_comb = 6'b000101;
 17'b00000000100001001 : data_comb = 6'b000110;
 17'b00000000100001010 : data_comb = 6'b001010;
 17'b00000000100001011 : data_comb = 6'b001010;
 17'b00000000100001100 : data_comb = 6'b001010;
 17'b00000000100001101 : data_comb = 6'b000101;
 17'b00000000100001110 : data_comb = 6'b000101;
 17'b00000000100001111 : data_comb = 6'b000101;
 17'b00000000100010000 : data_comb = 6'b000101;
 17'b00000000100010001 : data_comb = 6'b000101;
 17'b00000000100010010 : data_comb = 6'b000101;
 17'b00000000100010011 : data_comb = 6'b000101;
 17'b00000000100010100 : data_comb = 6'b000101;
 17'b00000000100010101 : data_comb = 6'b000101;
 17'b00000000100010110 : data_comb = 6'b000101;
 17'b00000000100010111 : data_comb = 6'b000101;
 17'b00000000100011000 : data_comb = 6'b000101;
 17'b00000000100011001 : data_comb = 6'b000101;
 17'b00000000100011010 : data_comb = 6'b000101;
 17'b00000000100011011 : data_comb = 6'b000101;
 17'b00000000100011100 : data_comb = 6'b000101;
 17'b00000000100011101 : data_comb = 6'b000101;
 17'b00000000100011110 : data_comb = 6'b000101;
 17'b00000000100011111 : data_comb = 6'b000101;
 17'b00000000100100000 : data_comb = 6'b000101;
 17'b00000000100100001 : data_comb = 6'b000101;
 17'b00000000100100010 : data_comb = 6'b000101;
 17'b00000000100100011 : data_comb = 6'b000101;
 17'b00000000100100100 : data_comb = 6'b000101;
 17'b00000000100100101 : data_comb = 6'b000101;
 17'b00000000100100110 : data_comb = 6'b000101;
 17'b00000000100100111 : data_comb = 6'b000101;
 17'b00000000100101000 : data_comb = 6'b000101;
 17'b00000000100101001 : data_comb = 6'b000101;
 17'b00000000100101010 : data_comb = 6'b000101;
 17'b00000000100101011 : data_comb = 6'b000101;
 17'b00000000100101100 : data_comb = 6'b000101;
 17'b00000000100101101 : data_comb = 6'b000101;
 17'b00000000100101110 : data_comb = 6'b000101;
 17'b00000000100101111 : data_comb = 6'b000101;
 17'b00000000100110000 : data_comb = 6'b000101;
 17'b00000000100110001 : data_comb = 6'b000101;
 17'b00000000100110010 : data_comb = 6'b000101;
 17'b00000000100110011 : data_comb = 6'b000101;
 17'b00000000100110100 : data_comb = 6'b000101;
 17'b00000000100110101 : data_comb = 6'b000101;
 17'b00000000100110110 : data_comb = 6'b000101;
 17'b00000000100110111 : data_comb = 6'b000101;
 17'b00000000100111000 : data_comb = 6'b000101;
 17'b00000000100111001 : data_comb = 6'b000101;
 17'b00000000100111010 : data_comb = 6'b000101;
 17'b00000000100111011 : data_comb = 6'b000101;
 17'b00000000100111100 : data_comb = 6'b000101;
 17'b00000000100111101 : data_comb = 6'b000101;
 17'b00000000100111110 : data_comb = 6'b000101;
 17'b00000000100111111 : data_comb = 6'b000101;
 17'b00000000101000000 : data_comb = 6'b000101;
 17'b00000000101000001 : data_comb = 6'b000101;
 17'b00000000101000010 : data_comb = 6'b000101;
 17'b00000000101000011 : data_comb = 6'b000101;
 17'b00000000101000100 : data_comb = 6'b000101;
 17'b00000000101000101 : data_comb = 6'b000101;
 17'b00000000101000110 : data_comb = 6'b000101;
 17'b00000000101000111 : data_comb = 6'b000101;
 17'b00000000101001000 : data_comb = 6'b000101;
 17'b00000000101001001 : data_comb = 6'b000101;
 17'b00000000101001010 : data_comb = 6'b101000;
 17'b00000000101001011 : data_comb = 6'b101000;
 17'b00000000101001100 : data_comb = 6'b111000;
 17'b00000000101001101 : data_comb = 6'b111000;
 17'b00000000101001110 : data_comb = 6'b111000;
 17'b00000000101001111 : data_comb = 6'b111000;
 17'b00000000101010000 : data_comb = 6'b010101;
 17'b00000000101010001 : data_comb = 6'b000101;
 17'b00000000101010010 : data_comb = 6'b000101;
 17'b00000000101010011 : data_comb = 6'b000101;
 17'b00000000101010100 : data_comb = 6'b000101;
 17'b00000000101010101 : data_comb = 6'b000101;
 17'b00000000101010110 : data_comb = 6'b000101;
 17'b00000000101010111 : data_comb = 6'b000110;
 17'b00000000101011000 : data_comb = 6'b000110;
 17'b00000000101011001 : data_comb = 6'b001010;
 17'b00000000101011010 : data_comb = 6'b001010;
 17'b00000000101011011 : data_comb = 6'b001010;
 17'b00000000101011100 : data_comb = 6'b001010;
 17'b00000000101011101 : data_comb = 6'b001010;
 17'b00000000101011110 : data_comb = 6'b000110;
 17'b00000000101011111 : data_comb = 6'b000101;
 17'b00000000101100000 : data_comb = 6'b000101;
 17'b00000000101100001 : data_comb = 6'b000101;
 17'b00000000101100010 : data_comb = 6'b000101;
 17'b00000000101100011 : data_comb = 6'b000101;
 17'b00000000101100100 : data_comb = 6'b000101;
 17'b00000000101100101 : data_comb = 6'b000101;
 17'b00000000101100110 : data_comb = 6'b000101;
 17'b00000000101100111 : data_comb = 6'b000101;
 17'b00000000101101000 : data_comb = 6'b000101;
 17'b00000000101101001 : data_comb = 6'b000101;
 17'b00000000101101010 : data_comb = 6'b000101;
 17'b00000000101101011 : data_comb = 6'b000101;
 17'b00000000101101100 : data_comb = 6'b000101;
 17'b00000000101101101 : data_comb = 6'b000101;
 17'b00000000101101110 : data_comb = 6'b000101;
 17'b00000000101101111 : data_comb = 6'b000101;
 17'b00000000101110000 : data_comb = 6'b000101;
 17'b00000000101110001 : data_comb = 6'b000101;
 17'b00000000101110010 : data_comb = 6'b000101;
 17'b00000000101110011 : data_comb = 6'b000101;
 17'b00000000101110100 : data_comb = 6'b000101;
 17'b00000000101110101 : data_comb = 6'b000101;
 17'b00000000101110110 : data_comb = 6'b000101;
 17'b00000000101110111 : data_comb = 6'b000101;
 17'b00000000101111000 : data_comb = 6'b000101;
 17'b00000000101111001 : data_comb = 6'b000101;
 17'b00000000101111010 : data_comb = 6'b000101;
 17'b00000000101111011 : data_comb = 6'b000101;
 17'b00000000101111100 : data_comb = 6'b000101;
 17'b00000000101111101 : data_comb = 6'b000101;
 17'b00000000101111110 : data_comb = 6'b000101;
 17'b00000000101111111 : data_comb = 6'b000101;
 17'b00000000110000000 : data_comb = 6'b000101;
 17'b00000000110000001 : data_comb = 6'b000101;
 17'b00000000110000010 : data_comb = 6'b000101;
 17'b00000000110000011 : data_comb = 6'b000101;
 17'b00000000110000100 : data_comb = 6'b000101;
 17'b00000000110000101 : data_comb = 6'b000101;
 17'b00000000110000110 : data_comb = 6'b000101;
 17'b00000000110000111 : data_comb = 6'b000101;
 17'b00000000110001000 : data_comb = 6'b000101;
 17'b00000000110001001 : data_comb = 6'b000101;
 17'b00000000110001010 : data_comb = 6'b000101;
 17'b00000000110001011 : data_comb = 6'b000101;
 17'b00000000110001100 : data_comb = 6'b000101;
 17'b00000000110001101 : data_comb = 6'b000101;
 17'b00000000110001110 : data_comb = 6'b000101;
 17'b00000000110001111 : data_comb = 6'b000101;
 17'b00000000110010000 : data_comb = 6'b000101;
 17'b00000000110010001 : data_comb = 6'b000101;
 17'b00000000110010010 : data_comb = 6'b000101;
 17'b00000000110010011 : data_comb = 6'b000101;
 17'b00000000110010100 : data_comb = 6'b000101;
 17'b00000000110010101 : data_comb = 6'b000101;
 17'b00000000110010110 : data_comb = 6'b000101;
 17'b00000000110010111 : data_comb = 6'b101000;
 17'b00000000110011000 : data_comb = 6'b101000;
 17'b00000000110011001 : data_comb = 6'b111000;
 17'b00000000110011010 : data_comb = 6'b111000;
 17'b00000000110011011 : data_comb = 6'b111000;
 17'b00000000110011100 : data_comb = 6'b111000;
 17'b00000000110011101 : data_comb = 6'b111000;
 17'b00000000110011110 : data_comb = 6'b111000;
 17'b00000000110011111 : data_comb = 6'b111000;
 17'b00000000110100000 : data_comb = 6'b010101;
 17'b00000000110100001 : data_comb = 6'b000101;
 17'b00000000110100010 : data_comb = 6'b000101;
 17'b00000000110100011 : data_comb = 6'b000101;
 17'b00000000110100100 : data_comb = 6'b000101;
 17'b00000000110100101 : data_comb = 6'b000101;
 17'b00000000110100110 : data_comb = 6'b000101;
 17'b00000000110100111 : data_comb = 6'b001010;
 17'b00000000110101000 : data_comb = 6'b001010;
 17'b00000000110101001 : data_comb = 6'b001010;
 17'b00000000110101010 : data_comb = 6'b001010;
 17'b00000000110101011 : data_comb = 6'b000110;
 17'b00000000110101100 : data_comb = 6'b000101;
 17'b00000000110101101 : data_comb = 6'b000101;
 17'b00000000110101110 : data_comb = 6'b000101;
 17'b00000000110101111 : data_comb = 6'b000101;
 17'b00000000110110000 : data_comb = 6'b000101;
 17'b00000000110110001 : data_comb = 6'b000101;
 17'b00000000110110010 : data_comb = 6'b000101;
 17'b00000000110110011 : data_comb = 6'b000101;
 17'b00000000110110100 : data_comb = 6'b000101;
 17'b00000000110110101 : data_comb = 6'b000101;
 17'b00000000110110110 : data_comb = 6'b000101;
 17'b00000000110110111 : data_comb = 6'b000101;
 17'b00000000110111000 : data_comb = 6'b000101;
 17'b00000000110111001 : data_comb = 6'b000101;
 17'b00000000110111010 : data_comb = 6'b000101;
 17'b00000000110111011 : data_comb = 6'b000101;
 17'b00000000110111100 : data_comb = 6'b000101;
 17'b00000000110111101 : data_comb = 6'b000101;
 17'b00000000110111110 : data_comb = 6'b000101;
 17'b00000000110111111 : data_comb = 6'b000101;
 17'b00000000111000000 : data_comb = 6'b000101;
 17'b00000000111000001 : data_comb = 6'b000101;
 17'b00000000111000010 : data_comb = 6'b000101;
 17'b00000000111000011 : data_comb = 6'b000101;
 17'b00000000111000100 : data_comb = 6'b000101;
 17'b00000000111000101 : data_comb = 6'b000101;
 17'b00000000111000110 : data_comb = 6'b000101;
 17'b00000000111000111 : data_comb = 6'b000101;
 17'b00000000111001000 : data_comb = 6'b000101;
 17'b00000000111001001 : data_comb = 6'b000101;
 17'b00000000111001010 : data_comb = 6'b101001;
 17'b00000000111001011 : data_comb = 6'b101000;
 17'b00000000111001100 : data_comb = 6'b010101;
 17'b00000000111001101 : data_comb = 6'b000101;
 17'b00000000111001110 : data_comb = 6'b000101;
 17'b00000000111001111 : data_comb = 6'b000101;
 17'b00000000111010000 : data_comb = 6'b000101;
 17'b00000000111010001 : data_comb = 6'b010101;
 17'b00000000111010010 : data_comb = 6'b010101;
 17'b00000000111010011 : data_comb = 6'b000101;
 17'b00000000111010100 : data_comb = 6'b000101;
 17'b00000000111010101 : data_comb = 6'b000101;
 17'b00000000111010110 : data_comb = 6'b000101;
 17'b00000000111010111 : data_comb = 6'b000101;
 17'b00000000111011000 : data_comb = 6'b000101;
 17'b00000000111011001 : data_comb = 6'b000101;
 17'b00000000111011010 : data_comb = 6'b000101;
 17'b00000000111011011 : data_comb = 6'b000101;
 17'b00000000111011100 : data_comb = 6'b000101;
 17'b00000000111011101 : data_comb = 6'b000101;
 17'b00000000111011110 : data_comb = 6'b000101;
 17'b00000000111011111 : data_comb = 6'b000101;
 17'b00000000111100000 : data_comb = 6'b000101;
 17'b00000000111100001 : data_comb = 6'b000101;
 17'b00000000111100010 : data_comb = 6'b000101;
 17'b00000000111100011 : data_comb = 6'b000101;
 17'b00000000111100100 : data_comb = 6'b000101;
 17'b00000000111100101 : data_comb = 6'b000101;
 17'b00000000111100110 : data_comb = 6'b000101;
 17'b00000000111100111 : data_comb = 6'b111000;
 17'b00000000111101000 : data_comb = 6'b111000;
 17'b00000000111101001 : data_comb = 6'b111000;
 17'b00000000111101010 : data_comb = 6'b111000;
 17'b00000000111101011 : data_comb = 6'b111000;
 17'b00000000111101100 : data_comb = 6'b111000;
 17'b00000000111101101 : data_comb = 6'b111000;
 17'b00000000111101110 : data_comb = 6'b111000;
 17'b00000000111101111 : data_comb = 6'b111000;
 17'b00000000111110000 : data_comb = 6'b101000;
 17'b00000000111110001 : data_comb = 6'b101000;
 17'b00000000111110010 : data_comb = 6'b000101;
 17'b00000000111110011 : data_comb = 6'b000101;
 17'b00000000111110100 : data_comb = 6'b000101;
 17'b00000000111110101 : data_comb = 6'b000101;
 17'b00000000111110110 : data_comb = 6'b001010;
 17'b00000000111110111 : data_comb = 6'b001010;
 17'b00000000111111000 : data_comb = 6'b001010;
 17'b00000000111111001 : data_comb = 6'b001010;
 17'b00000000111111010 : data_comb = 6'b000101;
 17'b00000000111111011 : data_comb = 6'b000101;
 17'b00000000111111100 : data_comb = 6'b000101;
 17'b00000000111111101 : data_comb = 6'b000101;
 17'b00000000111111110 : data_comb = 6'b000101;
 17'b00000000111111111 : data_comb = 6'b000101;
 17'b00000001000000000 : data_comb = 6'b000101;
 17'b00000001000000001 : data_comb = 6'b000101;
 17'b00000001000000010 : data_comb = 6'b000101;
 17'b00000001000000011 : data_comb = 6'b000101;
 17'b00000001000000100 : data_comb = 6'b000101;
 17'b00000001000000101 : data_comb = 6'b000101;
 17'b00000001000000110 : data_comb = 6'b000101;
 17'b00000001000000111 : data_comb = 6'b000101;
 17'b00000001000001000 : data_comb = 6'b000101;
 17'b00000001000001001 : data_comb = 6'b000101;
 17'b00000001000001010 : data_comb = 6'b000101;
 17'b00000001000001011 : data_comb = 6'b000101;
 17'b00000001000001100 : data_comb = 6'b000101;
 17'b00000001000001101 : data_comb = 6'b000101;
 17'b00000001000001110 : data_comb = 6'b000101;
 17'b00000001000001111 : data_comb = 6'b000101;
 17'b00000001000010000 : data_comb = 6'b000101;
 17'b00000001000010001 : data_comb = 6'b000101;
 17'b00000001000010010 : data_comb = 6'b000101;
 17'b00000001000010011 : data_comb = 6'b000101;
 17'b00000001000010100 : data_comb = 6'b000101;
 17'b00000001000010101 : data_comb = 6'b000101;
 17'b00000001000010110 : data_comb = 6'b000101;
 17'b00000001000010111 : data_comb = 6'b000101;
 17'b00000001000011000 : data_comb = 6'b010101;
 17'b00000001000011001 : data_comb = 6'b111000;
 17'b00000001000011010 : data_comb = 6'b111000;
 17'b00000001000011011 : data_comb = 6'b111000;
 17'b00000001000011100 : data_comb = 6'b111000;
 17'b00000001000011101 : data_comb = 6'b000101;
 17'b00000001000011110 : data_comb = 6'b000101;
 17'b00000001000011111 : data_comb = 6'b000101;
 17'b00000001000100000 : data_comb = 6'b101000;
 17'b00000001000100001 : data_comb = 6'b111000;
 17'b00000001000100010 : data_comb = 6'b111000;
 17'b00000001000100011 : data_comb = 6'b101000;
 17'b00000001000100100 : data_comb = 6'b000101;
 17'b00000001000100101 : data_comb = 6'b000101;
 17'b00000001000100110 : data_comb = 6'b000101;
 17'b00000001000100111 : data_comb = 6'b000101;
 17'b00000001000101000 : data_comb = 6'b000101;
 17'b00000001000101001 : data_comb = 6'b000101;
 17'b00000001000101010 : data_comb = 6'b000101;
 17'b00000001000101011 : data_comb = 6'b000101;
 17'b00000001000101100 : data_comb = 6'b000101;
 17'b00000001000101101 : data_comb = 6'b000101;
 17'b00000001000101110 : data_comb = 6'b000101;
 17'b00000001000101111 : data_comb = 6'b000101;
 17'b00000001000110000 : data_comb = 6'b000101;
 17'b00000001000110001 : data_comb = 6'b000101;
 17'b00000001000110010 : data_comb = 6'b000101;
 17'b00000001000110011 : data_comb = 6'b000101;
 17'b00000001000110100 : data_comb = 6'b000101;
 17'b00000001000110101 : data_comb = 6'b000101;
 17'b00000001000110110 : data_comb = 6'b000101;
 17'b00000001000110111 : data_comb = 6'b000101;
 17'b00000001000111000 : data_comb = 6'b000101;
 17'b00000001000111001 : data_comb = 6'b000101;
 17'b00000001000111010 : data_comb = 6'b010101;
 17'b00000001000111011 : data_comb = 6'b111000;
 17'b00000001000111100 : data_comb = 6'b111000;
 17'b00000001000111101 : data_comb = 6'b111000;
 17'b00000001000111110 : data_comb = 6'b111000;
 17'b00000001000111111 : data_comb = 6'b101000;
 17'b00000001001000000 : data_comb = 6'b101000;
 17'b00000001001000001 : data_comb = 6'b101000;
 17'b00000001001000010 : data_comb = 6'b000101;
 17'b00000001001000011 : data_comb = 6'b000101;
 17'b00000001001000100 : data_comb = 6'b000101;
 17'b00000001001000101 : data_comb = 6'b000110;
 17'b00000001001000110 : data_comb = 6'b001010;
 17'b00000001001000111 : data_comb = 6'b001010;
 17'b00000001001001000 : data_comb = 6'b001010;
 17'b00000001001001001 : data_comb = 6'b000110;
 17'b00000001001001010 : data_comb = 6'b000101;
 17'b00000001001001011 : data_comb = 6'b000101;
 17'b00000001001001100 : data_comb = 6'b000101;
 17'b00000001001001101 : data_comb = 6'b000101;
 17'b00000001001001110 : data_comb = 6'b000101;
 17'b00000001001001111 : data_comb = 6'b000101;
 17'b00000001001010000 : data_comb = 6'b000101;
 17'b00000001001010001 : data_comb = 6'b000101;
 17'b00000001001010010 : data_comb = 6'b000101;
 17'b00000001001010011 : data_comb = 6'b000101;
 17'b00000001001010100 : data_comb = 6'b000101;
 17'b00000001001010101 : data_comb = 6'b000101;
 17'b00000001001010110 : data_comb = 6'b000101;
 17'b00000001001010111 : data_comb = 6'b000101;
 17'b00000001001011000 : data_comb = 6'b000101;
 17'b00000001001011001 : data_comb = 6'b000101;
 17'b00000001001011010 : data_comb = 6'b000101;
 17'b00000001001011011 : data_comb = 6'b000101;
 17'b00000001001011100 : data_comb = 6'b000101;
 17'b00000001001011101 : data_comb = 6'b000101;
 17'b00000001001011110 : data_comb = 6'b000101;
 17'b00000001001011111 : data_comb = 6'b000101;
 17'b00000001001100000 : data_comb = 6'b000101;
 17'b00000001001100001 : data_comb = 6'b000101;
 17'b00000001001100010 : data_comb = 6'b000101;
 17'b00000001001100011 : data_comb = 6'b000101;
 17'b00000001001100100 : data_comb = 6'b000101;
 17'b00000001001100101 : data_comb = 6'b000101;
 17'b00000001001100110 : data_comb = 6'b000101;
 17'b00000001001100111 : data_comb = 6'b000101;
 17'b00000001001101000 : data_comb = 6'b101000;
 17'b00000001001101001 : data_comb = 6'b111000;
 17'b00000001001101010 : data_comb = 6'b111000;
 17'b00000001001101011 : data_comb = 6'b111000;
 17'b00000001001101100 : data_comb = 6'b111000;
 17'b00000001001101101 : data_comb = 6'b111000;
 17'b00000001001101110 : data_comb = 6'b000101;
 17'b00000001001101111 : data_comb = 6'b010101;
 17'b00000001001110000 : data_comb = 6'b111000;
 17'b00000001001110001 : data_comb = 6'b111000;
 17'b00000001001110010 : data_comb = 6'b111000;
 17'b00000001001110011 : data_comb = 6'b111000;
 17'b00000001001110100 : data_comb = 6'b010101;
 17'b00000001001110101 : data_comb = 6'b000101;
 17'b00000001001110110 : data_comb = 6'b000101;
 17'b00000001001110111 : data_comb = 6'b000101;
 17'b00000001001111000 : data_comb = 6'b000101;
 17'b00000001001111001 : data_comb = 6'b000101;
 17'b00000001001111010 : data_comb = 6'b000101;
 17'b00000001001111011 : data_comb = 6'b000101;
 17'b00000001001111100 : data_comb = 6'b000101;
 17'b00000001001111101 : data_comb = 6'b000101;
 17'b00000001001111110 : data_comb = 6'b000101;
 17'b00000001001111111 : data_comb = 6'b000101;
 17'b00000001010000000 : data_comb = 6'b000101;
 17'b00000001010000001 : data_comb = 6'b000101;
 17'b00000001010000010 : data_comb = 6'b000101;
 17'b00000001010000011 : data_comb = 6'b000101;
 17'b00000001010000100 : data_comb = 6'b000101;
 17'b00000001010000101 : data_comb = 6'b000101;
 17'b00000001010000110 : data_comb = 6'b000101;
 17'b00000001010000111 : data_comb = 6'b000101;
 17'b00000001010001000 : data_comb = 6'b000101;
 17'b00000001010001001 : data_comb = 6'b000101;
 17'b00000001010001010 : data_comb = 6'b000101;
 17'b00000001010001011 : data_comb = 6'b010101;
 17'b00000001010001100 : data_comb = 6'b010101;
 17'b00000001010001101 : data_comb = 6'b010101;
 17'b00000001010001110 : data_comb = 6'b010101;
 17'b00000001010001111 : data_comb = 6'b000101;
 17'b00000001010010000 : data_comb = 6'b000101;
 17'b00000001010010001 : data_comb = 6'b000101;
 17'b00000001010010010 : data_comb = 6'b000101;
 17'b00000001010010011 : data_comb = 6'b000101;
 17'b00000001010010100 : data_comb = 6'b000101;
 17'b00000001010010101 : data_comb = 6'b001010;
 17'b00000001010010110 : data_comb = 6'b001010;
 17'b00000001010010111 : data_comb = 6'b001010;
 17'b00000001010011000 : data_comb = 6'b001010;
 17'b00000001010011001 : data_comb = 6'b000110;
 17'b00000001010011010 : data_comb = 6'b000101;
 17'b00000001010011011 : data_comb = 6'b000101;
 17'b00000001010011100 : data_comb = 6'b000101;
 17'b00000001010011101 : data_comb = 6'b000101;
 17'b00000001010011110 : data_comb = 6'b000101;
 17'b00000001010011111 : data_comb = 6'b000101;
 17'b00000001010100000 : data_comb = 6'b000101;
 17'b00000001010100001 : data_comb = 6'b000101;
 17'b00000001010100010 : data_comb = 6'b000101;
 17'b00000001010100011 : data_comb = 6'b000101;
 17'b00000001010100100 : data_comb = 6'b000101;
 17'b00000001010100101 : data_comb = 6'b000101;
 17'b00000001010100110 : data_comb = 6'b000101;
 17'b00000001010100111 : data_comb = 6'b000101;
 17'b00000001010101000 : data_comb = 6'b000101;
 17'b00000001010101001 : data_comb = 6'b000101;
 17'b00000001010101010 : data_comb = 6'b000101;
 17'b00000001010101011 : data_comb = 6'b000101;
 17'b00000001010101100 : data_comb = 6'b000101;
 17'b00000001010101101 : data_comb = 6'b000101;
 17'b00000001010101110 : data_comb = 6'b000101;
 17'b00000001010101111 : data_comb = 6'b000101;
 17'b00000001010110000 : data_comb = 6'b000101;
 17'b00000001010110001 : data_comb = 6'b000101;
 17'b00000001010110010 : data_comb = 6'b000101;
 17'b00000001010110011 : data_comb = 6'b000101;
 17'b00000001010110100 : data_comb = 6'b000101;
 17'b00000001010110101 : data_comb = 6'b000101;
 17'b00000001010110110 : data_comb = 6'b000101;
 17'b00000001010110111 : data_comb = 6'b011001;
 17'b00000001010111000 : data_comb = 6'b111000;
 17'b00000001010111001 : data_comb = 6'b111000;
 17'b00000001010111010 : data_comb = 6'b111000;
 17'b00000001010111011 : data_comb = 6'b111000;
 17'b00000001010111100 : data_comb = 6'b111000;
 17'b00000001010111101 : data_comb = 6'b111000;
 17'b00000001010111110 : data_comb = 6'b111000;
 17'b00000001010111111 : data_comb = 6'b111000;
 17'b00000001011000000 : data_comb = 6'b111000;
 17'b00000001011000001 : data_comb = 6'b111000;
 17'b00000001011000010 : data_comb = 6'b111000;
 17'b00000001011000011 : data_comb = 6'b111000;
 17'b00000001011000100 : data_comb = 6'b000101;
 17'b00000001011000101 : data_comb = 6'b000101;
 17'b00000001011000110 : data_comb = 6'b000101;
 17'b00000001011000111 : data_comb = 6'b000101;
 17'b00000001011001000 : data_comb = 6'b101000;
 17'b00000001011001001 : data_comb = 6'b101000;
 17'b00000001011001010 : data_comb = 6'b101000;
 17'b00000001011001011 : data_comb = 6'b000101;
 17'b00000001011001100 : data_comb = 6'b000101;
 17'b00000001011001101 : data_comb = 6'b000101;
 17'b00000001011001110 : data_comb = 6'b000101;
 17'b00000001011001111 : data_comb = 6'b000101;
 17'b00000001011010000 : data_comb = 6'b000101;
 17'b00000001011010001 : data_comb = 6'b000101;
 17'b00000001011010010 : data_comb = 6'b000101;
 17'b00000001011010011 : data_comb = 6'b000101;
 17'b00000001011010100 : data_comb = 6'b000101;
 17'b00000001011010101 : data_comb = 6'b000101;
 17'b00000001011010110 : data_comb = 6'b000101;
 17'b00000001011010111 : data_comb = 6'b000101;
 17'b00000001011011000 : data_comb = 6'b000101;
 17'b00000001011011001 : data_comb = 6'b000101;
 17'b00000001011011010 : data_comb = 6'b000101;
 17'b00000001011011011 : data_comb = 6'b000101;
 17'b00000001011011100 : data_comb = 6'b000101;
 17'b00000001011011101 : data_comb = 6'b000101;
 17'b00000001011011110 : data_comb = 6'b000101;
 17'b00000001011011111 : data_comb = 6'b000101;
 17'b00000001011100000 : data_comb = 6'b000101;
 17'b00000001011100001 : data_comb = 6'b000101;
 17'b00000001011100010 : data_comb = 6'b000101;
 17'b00000001011100011 : data_comb = 6'b000101;
 17'b00000001011100100 : data_comb = 6'b000110;
 17'b00000001011100101 : data_comb = 6'b001010;
 17'b00000001011100110 : data_comb = 6'b001010;
 17'b00000001011100111 : data_comb = 6'b001010;
 17'b00000001011101000 : data_comb = 6'b000110;
 17'b00000001011101001 : data_comb = 6'b000101;
 17'b00000001011101010 : data_comb = 6'b000101;
 17'b00000001011101011 : data_comb = 6'b000101;
 17'b00000001011101100 : data_comb = 6'b000101;
 17'b00000001011101101 : data_comb = 6'b000101;
 17'b00000001011101110 : data_comb = 6'b000101;
 17'b00000001011101111 : data_comb = 6'b000101;
 17'b00000001011110000 : data_comb = 6'b000101;
 17'b00000001011110001 : data_comb = 6'b000101;
 17'b00000001011110010 : data_comb = 6'b000101;
 17'b00000001011110011 : data_comb = 6'b000101;
 17'b00000001011110100 : data_comb = 6'b000101;
 17'b00000001011110101 : data_comb = 6'b000101;
 17'b00000001011110110 : data_comb = 6'b000101;
 17'b00000001011110111 : data_comb = 6'b000101;
 17'b00000001011111000 : data_comb = 6'b000101;
 17'b00000001011111001 : data_comb = 6'b000101;
 17'b00000001011111010 : data_comb = 6'b000101;
 17'b00000001011111011 : data_comb = 6'b000101;
 17'b00000001011111100 : data_comb = 6'b000101;
 17'b00000001011111101 : data_comb = 6'b000101;
 17'b00000001011111110 : data_comb = 6'b000101;
 17'b00000001011111111 : data_comb = 6'b000101;
 17'b00000001100000000 : data_comb = 6'b000101;
 17'b00000001100000001 : data_comb = 6'b000101;
 17'b00000001100000010 : data_comb = 6'b000101;
 17'b00000001100000011 : data_comb = 6'b000101;
 17'b00000001100000100 : data_comb = 6'b000101;
 17'b00000001100000101 : data_comb = 6'b000101;
 17'b00000001100000110 : data_comb = 6'b000101;
 17'b00000001100000111 : data_comb = 6'b011001;
 17'b00000001100001000 : data_comb = 6'b111000;
 17'b00000001100001001 : data_comb = 6'b111000;
 17'b00000001100001010 : data_comb = 6'b111000;
 17'b00000001100001011 : data_comb = 6'b111000;
 17'b00000001100001100 : data_comb = 6'b111000;
 17'b00000001100001101 : data_comb = 6'b111000;
 17'b00000001100001110 : data_comb = 6'b111000;
 17'b00000001100001111 : data_comb = 6'b111000;
 17'b00000001100010000 : data_comb = 6'b111000;
 17'b00000001100010001 : data_comb = 6'b111000;
 17'b00000001100010010 : data_comb = 6'b111000;
 17'b00000001100010011 : data_comb = 6'b101000;
 17'b00000001100010100 : data_comb = 6'b000101;
 17'b00000001100010101 : data_comb = 6'b000101;
 17'b00000001100010110 : data_comb = 6'b000101;
 17'b00000001100010111 : data_comb = 6'b101000;
 17'b00000001100011000 : data_comb = 6'b111000;
 17'b00000001100011001 : data_comb = 6'b111000;
 17'b00000001100011010 : data_comb = 6'b111000;
 17'b00000001100011011 : data_comb = 6'b111000;
 17'b00000001100011100 : data_comb = 6'b000101;
 17'b00000001100011101 : data_comb = 6'b000101;
 17'b00000001100011110 : data_comb = 6'b000101;
 17'b00000001100011111 : data_comb = 6'b000101;
 17'b00000001100100000 : data_comb = 6'b000101;
 17'b00000001100100001 : data_comb = 6'b000101;
 17'b00000001100100010 : data_comb = 6'b000101;
 17'b00000001100100011 : data_comb = 6'b000101;
 17'b00000001100100100 : data_comb = 6'b000101;
 17'b00000001100100101 : data_comb = 6'b101000;
 17'b00000001100100110 : data_comb = 6'b101000;
 17'b00000001100100111 : data_comb = 6'b010101;
 17'b00000001100101000 : data_comb = 6'b000101;
 17'b00000001100101001 : data_comb = 6'b000101;
 17'b00000001100101010 : data_comb = 6'b000101;
 17'b00000001100101011 : data_comb = 6'b000101;
 17'b00000001100101100 : data_comb = 6'b000101;
 17'b00000001100101101 : data_comb = 6'b000101;
 17'b00000001100101110 : data_comb = 6'b000101;
 17'b00000001100101111 : data_comb = 6'b000101;
 17'b00000001100110000 : data_comb = 6'b000101;
 17'b00000001100110001 : data_comb = 6'b000101;
 17'b00000001100110010 : data_comb = 6'b000101;
 17'b00000001100110011 : data_comb = 6'b000101;
 17'b00000001100110100 : data_comb = 6'b000110;
 17'b00000001100110101 : data_comb = 6'b001010;
 17'b00000001100110110 : data_comb = 6'b001010;
 17'b00000001100110111 : data_comb = 6'b001010;
 17'b00000001100111000 : data_comb = 6'b000110;
 17'b00000001100111001 : data_comb = 6'b000101;
 17'b00000001100111010 : data_comb = 6'b000101;
 17'b00000001100111011 : data_comb = 6'b000101;
 17'b00000001100111100 : data_comb = 6'b000101;
 17'b00000001100111101 : data_comb = 6'b000101;
 17'b00000001100111110 : data_comb = 6'b000101;
 17'b00000001100111111 : data_comb = 6'b000101;
 17'b00000001101000000 : data_comb = 6'b000101;
 17'b00000001101000001 : data_comb = 6'b000101;
 17'b00000001101000010 : data_comb = 6'b000101;
 17'b00000001101000011 : data_comb = 6'b000101;
 17'b00000001101000100 : data_comb = 6'b000101;
 17'b00000001101000101 : data_comb = 6'b000101;
 17'b00000001101000110 : data_comb = 6'b000101;
 17'b00000001101000111 : data_comb = 6'b000101;
 17'b00000001101001000 : data_comb = 6'b000101;
 17'b00000001101001001 : data_comb = 6'b000101;
 17'b00000001101001010 : data_comb = 6'b000101;
 17'b00000001101001011 : data_comb = 6'b000101;
 17'b00000001101001100 : data_comb = 6'b000101;
 17'b00000001101001101 : data_comb = 6'b000101;
 17'b00000001101001110 : data_comb = 6'b000101;
 17'b00000001101001111 : data_comb = 6'b000101;
 17'b00000001101010000 : data_comb = 6'b000101;
 17'b00000001101010001 : data_comb = 6'b000101;
 17'b00000001101010010 : data_comb = 6'b000101;
 17'b00000001101010011 : data_comb = 6'b000101;
 17'b00000001101010100 : data_comb = 6'b000101;
 17'b00000001101010101 : data_comb = 6'b000101;
 17'b00000001101010110 : data_comb = 6'b000101;
 17'b00000001101010111 : data_comb = 6'b011001;
 17'b00000001101011000 : data_comb = 6'b111000;
 17'b00000001101011001 : data_comb = 6'b111000;
 17'b00000001101011010 : data_comb = 6'b111000;
 17'b00000001101011011 : data_comb = 6'b111000;
 17'b00000001101011100 : data_comb = 6'b111000;
 17'b00000001101011101 : data_comb = 6'b111000;
 17'b00000001101011110 : data_comb = 6'b111000;
 17'b00000001101011111 : data_comb = 6'b111000;
 17'b00000001101100000 : data_comb = 6'b111000;
 17'b00000001101100001 : data_comb = 6'b101000;
 17'b00000001101100010 : data_comb = 6'b000101;
 17'b00000001101100011 : data_comb = 6'b000101;
 17'b00000001101100100 : data_comb = 6'b000101;
 17'b00000001101100101 : data_comb = 6'b000101;
 17'b00000001101100110 : data_comb = 6'b111000;
 17'b00000001101100111 : data_comb = 6'b111000;
 17'b00000001101101000 : data_comb = 6'b111000;
 17'b00000001101101001 : data_comb = 6'b111000;
 17'b00000001101101010 : data_comb = 6'b111000;
 17'b00000001101101011 : data_comb = 6'b111000;
 17'b00000001101101100 : data_comb = 6'b101000;
 17'b00000001101101101 : data_comb = 6'b000101;
 17'b00000001101101110 : data_comb = 6'b000101;
 17'b00000001101101111 : data_comb = 6'b000101;
 17'b00000001101110000 : data_comb = 6'b000101;
 17'b00000001101110001 : data_comb = 6'b000101;
 17'b00000001101110010 : data_comb = 6'b000101;
 17'b00000001101110011 : data_comb = 6'b010101;
 17'b00000001101110100 : data_comb = 6'b111000;
 17'b00000001101110101 : data_comb = 6'b111000;
 17'b00000001101110110 : data_comb = 6'b111000;
 17'b00000001101110111 : data_comb = 6'b111000;
 17'b00000001101111000 : data_comb = 6'b111000;
 17'b00000001101111001 : data_comb = 6'b000101;
 17'b00000001101111010 : data_comb = 6'b000101;
 17'b00000001101111011 : data_comb = 6'b000101;
 17'b00000001101111100 : data_comb = 6'b000101;
 17'b00000001101111101 : data_comb = 6'b000101;
 17'b00000001101111110 : data_comb = 6'b000101;
 17'b00000001101111111 : data_comb = 6'b000101;
 17'b00000001110000000 : data_comb = 6'b000101;
 17'b00000001110000001 : data_comb = 6'b000101;
 17'b00000001110000010 : data_comb = 6'b000101;
 17'b00000001110000011 : data_comb = 6'b000101;
 17'b00000001110000100 : data_comb = 6'b000110;
 17'b00000001110000101 : data_comb = 6'b001010;
 17'b00000001110000110 : data_comb = 6'b001010;
 17'b00000001110000111 : data_comb = 6'b001010;
 17'b00000001110001000 : data_comb = 6'b000110;
 17'b00000001110001001 : data_comb = 6'b000101;
 17'b00000001110001010 : data_comb = 6'b000101;
 17'b00000001110001011 : data_comb = 6'b000101;
 17'b00000001110001100 : data_comb = 6'b000101;
 17'b00000001110001101 : data_comb = 6'b000101;
 17'b00000001110001110 : data_comb = 6'b000101;
 17'b00000001110001111 : data_comb = 6'b000101;
 17'b00000001110010000 : data_comb = 6'b000101;
 17'b00000001110010001 : data_comb = 6'b000101;
 17'b00000001110010010 : data_comb = 6'b000101;
 17'b00000001110010011 : data_comb = 6'b000101;
 17'b00000001110010100 : data_comb = 6'b000101;
 17'b00000001110010101 : data_comb = 6'b000101;
 17'b00000001110010110 : data_comb = 6'b000101;
 17'b00000001110010111 : data_comb = 6'b111000;
 17'b00000001110011000 : data_comb = 6'b111000;
 17'b00000001110011001 : data_comb = 6'b101001;
 17'b00000001110011010 : data_comb = 6'b000101;
 17'b00000001110011011 : data_comb = 6'b000101;
 17'b00000001110011100 : data_comb = 6'b000101;
 17'b00000001110011101 : data_comb = 6'b000101;
 17'b00000001110011110 : data_comb = 6'b000101;
 17'b00000001110011111 : data_comb = 6'b000101;
 17'b00000001110100000 : data_comb = 6'b000101;
 17'b00000001110100001 : data_comb = 6'b000101;
 17'b00000001110100010 : data_comb = 6'b000101;
 17'b00000001110100011 : data_comb = 6'b000101;
 17'b00000001110100100 : data_comb = 6'b000101;
 17'b00000001110100101 : data_comb = 6'b000101;
 17'b00000001110100110 : data_comb = 6'b000101;
 17'b00000001110100111 : data_comb = 6'b000101;
 17'b00000001110101000 : data_comb = 6'b101000;
 17'b00000001110101001 : data_comb = 6'b111000;
 17'b00000001110101010 : data_comb = 6'b111000;
 17'b00000001110101011 : data_comb = 6'b111000;
 17'b00000001110101100 : data_comb = 6'b111000;
 17'b00000001110101101 : data_comb = 6'b111000;
 17'b00000001110101110 : data_comb = 6'b111000;
 17'b00000001110101111 : data_comb = 6'b111000;
 17'b00000001110110000 : data_comb = 6'b111000;
 17'b00000001110110001 : data_comb = 6'b000101;
 17'b00000001110110010 : data_comb = 6'b000101;
 17'b00000001110110011 : data_comb = 6'b000101;
 17'b00000001110110100 : data_comb = 6'b000101;
 17'b00000001110110101 : data_comb = 6'b010101;
 17'b00000001110110110 : data_comb = 6'b101000;
 17'b00000001110110111 : data_comb = 6'b101000;
 17'b00000001110111000 : data_comb = 6'b101000;
 17'b00000001110111001 : data_comb = 6'b101001;
 17'b00000001110111010 : data_comb = 6'b101000;
 17'b00000001110111011 : data_comb = 6'b101000;
 17'b00000001110111100 : data_comb = 6'b101000;
 17'b00000001110111101 : data_comb = 6'b000101;
 17'b00000001110111110 : data_comb = 6'b000101;
 17'b00000001110111111 : data_comb = 6'b000101;
 17'b00000001111000000 : data_comb = 6'b111000;
 17'b00000001111000001 : data_comb = 6'b101000;
 17'b00000001111000010 : data_comb = 6'b010101;
 17'b00000001111000011 : data_comb = 6'b101000;
 17'b00000001111000100 : data_comb = 6'b111000;
 17'b00000001111000101 : data_comb = 6'b111000;
 17'b00000001111000110 : data_comb = 6'b111000;
 17'b00000001111000111 : data_comb = 6'b111000;
 17'b00000001111001000 : data_comb = 6'b111000;
 17'b00000001111001001 : data_comb = 6'b010101;
 17'b00000001111001010 : data_comb = 6'b000101;
 17'b00000001111001011 : data_comb = 6'b000101;
 17'b00000001111001100 : data_comb = 6'b000101;
 17'b00000001111001101 : data_comb = 6'b000101;
 17'b00000001111001110 : data_comb = 6'b000101;
 17'b00000001111001111 : data_comb = 6'b000101;
 17'b00000001111010000 : data_comb = 6'b000101;
 17'b00000001111010001 : data_comb = 6'b000101;
 17'b00000001111010010 : data_comb = 6'b000101;
 17'b00000001111010011 : data_comb = 6'b000101;
 17'b00000001111010100 : data_comb = 6'b000110;
 17'b00000001111010101 : data_comb = 6'b001010;
 17'b00000001111010110 : data_comb = 6'b001010;
 17'b00000001111010111 : data_comb = 6'b001010;
 17'b00000001111011000 : data_comb = 6'b000110;
 17'b00000001111011001 : data_comb = 6'b000101;
 17'b00000001111011010 : data_comb = 6'b000101;
 17'b00000001111011011 : data_comb = 6'b000101;
 17'b00000001111011100 : data_comb = 6'b000101;
 17'b00000001111011101 : data_comb = 6'b000101;
 17'b00000001111011110 : data_comb = 6'b000101;
 17'b00000001111011111 : data_comb = 6'b000101;
 17'b00000001111100000 : data_comb = 6'b000101;
 17'b00000001111100001 : data_comb = 6'b000101;
 17'b00000001111100010 : data_comb = 6'b000101;
 17'b00000001111100011 : data_comb = 6'b000101;
 17'b00000001111100100 : data_comb = 6'b000101;
 17'b00000001111100101 : data_comb = 6'b000101;
 17'b00000001111100110 : data_comb = 6'b101000;
 17'b00000001111100111 : data_comb = 6'b111000;
 17'b00000001111101000 : data_comb = 6'b111000;
 17'b00000001111101001 : data_comb = 6'b111000;
 17'b00000001111101010 : data_comb = 6'b000101;
 17'b00000001111101011 : data_comb = 6'b000101;
 17'b00000001111101100 : data_comb = 6'b000101;
 17'b00000001111101101 : data_comb = 6'b000101;
 17'b00000001111101110 : data_comb = 6'b000101;
 17'b00000001111101111 : data_comb = 6'b000101;
 17'b00000001111110000 : data_comb = 6'b000101;
 17'b00000001111110001 : data_comb = 6'b000101;
 17'b00000001111110010 : data_comb = 6'b000101;
 17'b00000001111110011 : data_comb = 6'b101000;
 17'b00000001111110100 : data_comb = 6'b101000;
 17'b00000001111110101 : data_comb = 6'b000101;
 17'b00000001111110110 : data_comb = 6'b000101;
 17'b00000001111110111 : data_comb = 6'b000101;
 17'b00000001111111000 : data_comb = 6'b111000;
 17'b00000001111111001 : data_comb = 6'b111000;
 17'b00000001111111010 : data_comb = 6'b111000;
 17'b00000001111111011 : data_comb = 6'b111000;
 17'b00000001111111100 : data_comb = 6'b111000;
 17'b00000001111111101 : data_comb = 6'b111000;
 17'b00000001111111110 : data_comb = 6'b111000;
 17'b00000001111111111 : data_comb = 6'b111000;
 17'b00000010000000000 : data_comb = 6'b111000;
 17'b00000010000000001 : data_comb = 6'b111000;
 17'b00000010000000010 : data_comb = 6'b101000;
 17'b00000010000000011 : data_comb = 6'b000101;
 17'b00000010000000100 : data_comb = 6'b000101;
 17'b00000010000000101 : data_comb = 6'b000101;
 17'b00000010000000110 : data_comb = 6'b000101;
 17'b00000010000000111 : data_comb = 6'b000101;
 17'b00000010000001000 : data_comb = 6'b000101;
 17'b00000010000001001 : data_comb = 6'b000101;
 17'b00000010000001010 : data_comb = 6'b000101;
 17'b00000010000001011 : data_comb = 6'b000101;
 17'b00000010000001100 : data_comb = 6'b000101;
 17'b00000010000001101 : data_comb = 6'b000101;
 17'b00000010000001110 : data_comb = 6'b000101;
 17'b00000010000001111 : data_comb = 6'b000101;
 17'b00000010000010000 : data_comb = 6'b111000;
 17'b00000010000010001 : data_comb = 6'b111000;
 17'b00000010000010010 : data_comb = 6'b111000;
 17'b00000010000010011 : data_comb = 6'b111000;
 17'b00000010000010100 : data_comb = 6'b111000;
 17'b00000010000010101 : data_comb = 6'b111000;
 17'b00000010000010110 : data_comb = 6'b111000;
 17'b00000010000010111 : data_comb = 6'b111000;
 17'b00000010000011000 : data_comb = 6'b111000;
 17'b00000010000011001 : data_comb = 6'b101001;
 17'b00000010000011010 : data_comb = 6'b000101;
 17'b00000010000011011 : data_comb = 6'b010101;
 17'b00000010000011100 : data_comb = 6'b111000;
 17'b00000010000011101 : data_comb = 6'b111000;
 17'b00000010000011110 : data_comb = 6'b000101;
 17'b00000010000011111 : data_comb = 6'b000101;
 17'b00000010000100000 : data_comb = 6'b000101;
 17'b00000010000100001 : data_comb = 6'b000101;
 17'b00000010000100010 : data_comb = 6'b000101;
 17'b00000010000100011 : data_comb = 6'b000101;
 17'b00000010000100100 : data_comb = 6'b000110;
 17'b00000010000100101 : data_comb = 6'b001010;
 17'b00000010000100110 : data_comb = 6'b001010;
 17'b00000010000100111 : data_comb = 6'b001010;
 17'b00000010000101000 : data_comb = 6'b001010;
 17'b00000010000101001 : data_comb = 6'b000101;
 17'b00000010000101010 : data_comb = 6'b000101;
 17'b00000010000101011 : data_comb = 6'b000101;
 17'b00000010000101100 : data_comb = 6'b000101;
 17'b00000010000101101 : data_comb = 6'b000101;
 17'b00000010000101110 : data_comb = 6'b000101;
 17'b00000010000101111 : data_comb = 6'b000101;
 17'b00000010000110000 : data_comb = 6'b000101;
 17'b00000010000110001 : data_comb = 6'b000101;
 17'b00000010000110010 : data_comb = 6'b000101;
 17'b00000010000110011 : data_comb = 6'b000101;
 17'b00000010000110100 : data_comb = 6'b111000;
 17'b00000010000110101 : data_comb = 6'b111000;
 17'b00000010000110110 : data_comb = 6'b111000;
 17'b00000010000110111 : data_comb = 6'b111000;
 17'b00000010000111000 : data_comb = 6'b111000;
 17'b00000010000111001 : data_comb = 6'b111000;
 17'b00000010000111010 : data_comb = 6'b111000;
 17'b00000010000111011 : data_comb = 6'b111000;
 17'b00000010000111100 : data_comb = 6'b010101;
 17'b00000010000111101 : data_comb = 6'b000101;
 17'b00000010000111110 : data_comb = 6'b000101;
 17'b00000010000111111 : data_comb = 6'b000101;
 17'b00000010001000000 : data_comb = 6'b000101;
 17'b00000010001000001 : data_comb = 6'b000101;
 17'b00000010001000010 : data_comb = 6'b101000;
 17'b00000010001000011 : data_comb = 6'b111000;
 17'b00000010001000100 : data_comb = 6'b111000;
 17'b00000010001000101 : data_comb = 6'b111000;
 17'b00000010001000110 : data_comb = 6'b111000;
 17'b00000010001000111 : data_comb = 6'b111000;
 17'b00000010001001000 : data_comb = 6'b111000;
 17'b00000010001001001 : data_comb = 6'b111000;
 17'b00000010001001010 : data_comb = 6'b111000;
 17'b00000010001001011 : data_comb = 6'b111000;
 17'b00000010001001100 : data_comb = 6'b111000;
 17'b00000010001001101 : data_comb = 6'b111000;
 17'b00000010001001110 : data_comb = 6'b111000;
 17'b00000010001001111 : data_comb = 6'b111000;
 17'b00000010001010000 : data_comb = 6'b100101;
 17'b00000010001010001 : data_comb = 6'b100101;
 17'b00000010001010010 : data_comb = 6'b010101;
 17'b00000010001010011 : data_comb = 6'b000101;
 17'b00000010001010100 : data_comb = 6'b000101;
 17'b00000010001010101 : data_comb = 6'b000101;
 17'b00000010001010110 : data_comb = 6'b000101;
 17'b00000010001010111 : data_comb = 6'b000101;
 17'b00000010001011000 : data_comb = 6'b000101;
 17'b00000010001011001 : data_comb = 6'b000101;
 17'b00000010001011010 : data_comb = 6'b000101;
 17'b00000010001011011 : data_comb = 6'b000101;
 17'b00000010001011100 : data_comb = 6'b000101;
 17'b00000010001011101 : data_comb = 6'b000101;
 17'b00000010001011110 : data_comb = 6'b000101;
 17'b00000010001011111 : data_comb = 6'b000101;
 17'b00000010001100000 : data_comb = 6'b111000;
 17'b00000010001100001 : data_comb = 6'b111000;
 17'b00000010001100010 : data_comb = 6'b111000;
 17'b00000010001100011 : data_comb = 6'b111000;
 17'b00000010001100100 : data_comb = 6'b111000;
 17'b00000010001100101 : data_comb = 6'b111000;
 17'b00000010001100110 : data_comb = 6'b111000;
 17'b00000010001100111 : data_comb = 6'b111000;
 17'b00000010001101000 : data_comb = 6'b111000;
 17'b00000010001101001 : data_comb = 6'b111000;
 17'b00000010001101010 : data_comb = 6'b101000;
 17'b00000010001101011 : data_comb = 6'b111000;
 17'b00000010001101100 : data_comb = 6'b111000;
 17'b00000010001101101 : data_comb = 6'b111000;
 17'b00000010001101110 : data_comb = 6'b111000;
 17'b00000010001101111 : data_comb = 6'b000101;
 17'b00000010001110000 : data_comb = 6'b000101;
 17'b00000010001110001 : data_comb = 6'b000101;
 17'b00000010001110010 : data_comb = 6'b000101;
 17'b00000010001110011 : data_comb = 6'b000101;
 17'b00000010001110100 : data_comb = 6'b000101;
 17'b00000010001110101 : data_comb = 6'b000110;
 17'b00000010001110110 : data_comb = 6'b001010;
 17'b00000010001110111 : data_comb = 6'b001010;
 17'b00000010001111000 : data_comb = 6'b001010;
 17'b00000010001111001 : data_comb = 6'b000110;
 17'b00000010001111010 : data_comb = 6'b000101;
 17'b00000010001111011 : data_comb = 6'b000101;
 17'b00000010001111100 : data_comb = 6'b000101;
 17'b00000010001111101 : data_comb = 6'b000101;
 17'b00000010001111110 : data_comb = 6'b000101;
 17'b00000010001111111 : data_comb = 6'b000101;
 17'b00000010010000000 : data_comb = 6'b000101;
 17'b00000010010000001 : data_comb = 6'b000101;
 17'b00000010010000010 : data_comb = 6'b000101;
 17'b00000010010000011 : data_comb = 6'b000101;
 17'b00000010010000100 : data_comb = 6'b000101;
 17'b00000010010000101 : data_comb = 6'b000101;
 17'b00000010010000110 : data_comb = 6'b000101;
 17'b00000010010000111 : data_comb = 6'b000101;
 17'b00000010010001000 : data_comb = 6'b000101;
 17'b00000010010001001 : data_comb = 6'b000101;
 17'b00000010010001010 : data_comb = 6'b000101;
 17'b00000010010001011 : data_comb = 6'b010101;
 17'b00000010010001100 : data_comb = 6'b000101;
 17'b00000010010001101 : data_comb = 6'b000101;
 17'b00000010010001110 : data_comb = 6'b000101;
 17'b00000010010001111 : data_comb = 6'b000101;
 17'b00000010010010000 : data_comb = 6'b000101;
 17'b00000010010010001 : data_comb = 6'b000101;
 17'b00000010010010010 : data_comb = 6'b111000;
 17'b00000010010010011 : data_comb = 6'b111000;
 17'b00000010010010100 : data_comb = 6'b111000;
 17'b00000010010010101 : data_comb = 6'b111000;
 17'b00000010010010110 : data_comb = 6'b111000;
 17'b00000010010010111 : data_comb = 6'b111000;
 17'b00000010010011000 : data_comb = 6'b111000;
 17'b00000010010011001 : data_comb = 6'b111000;
 17'b00000010010011010 : data_comb = 6'b111000;
 17'b00000010010011011 : data_comb = 6'b111000;
 17'b00000010010011100 : data_comb = 6'b111000;
 17'b00000010010011101 : data_comb = 6'b000101;
 17'b00000010010011110 : data_comb = 6'b000101;
 17'b00000010010011111 : data_comb = 6'b000101;
 17'b00000010010100000 : data_comb = 6'b000101;
 17'b00000010010100001 : data_comb = 6'b000101;
 17'b00000010010100010 : data_comb = 6'b000101;
 17'b00000010010100011 : data_comb = 6'b000101;
 17'b00000010010100100 : data_comb = 6'b000101;
 17'b00000010010100101 : data_comb = 6'b000101;
 17'b00000010010100110 : data_comb = 6'b000101;
 17'b00000010010100111 : data_comb = 6'b000101;
 17'b00000010010101000 : data_comb = 6'b000101;
 17'b00000010010101001 : data_comb = 6'b000101;
 17'b00000010010101010 : data_comb = 6'b000101;
 17'b00000010010101011 : data_comb = 6'b000101;
 17'b00000010010101100 : data_comb = 6'b000101;
 17'b00000010010101101 : data_comb = 6'b000101;
 17'b00000010010101110 : data_comb = 6'b000101;
 17'b00000010010101111 : data_comb = 6'b000101;
 17'b00000010010110000 : data_comb = 6'b111000;
 17'b00000010010110001 : data_comb = 6'b111000;
 17'b00000010010110010 : data_comb = 6'b111000;
 17'b00000010010110011 : data_comb = 6'b111000;
 17'b00000010010110100 : data_comb = 6'b111000;
 17'b00000010010110101 : data_comb = 6'b111000;
 17'b00000010010110110 : data_comb = 6'b111000;
 17'b00000010010110111 : data_comb = 6'b111000;
 17'b00000010010111000 : data_comb = 6'b111000;
 17'b00000010010111001 : data_comb = 6'b111000;
 17'b00000010010111010 : data_comb = 6'b111000;
 17'b00000010010111011 : data_comb = 6'b111000;
 17'b00000010010111100 : data_comb = 6'b111000;
 17'b00000010010111101 : data_comb = 6'b111000;
 17'b00000010010111110 : data_comb = 6'b111000;
 17'b00000010010111111 : data_comb = 6'b000101;
 17'b00000010011000000 : data_comb = 6'b000101;
 17'b00000010011000001 : data_comb = 6'b000101;
 17'b00000010011000010 : data_comb = 6'b000101;
 17'b00000010011000011 : data_comb = 6'b000101;
 17'b00000010011000100 : data_comb = 6'b000101;
 17'b00000010011000101 : data_comb = 6'b000110;
 17'b00000010011000110 : data_comb = 6'b001010;
 17'b00000010011000111 : data_comb = 6'b001010;
 17'b00000010011001000 : data_comb = 6'b001010;
 17'b00000010011001001 : data_comb = 6'b001010;
 17'b00000010011001010 : data_comb = 6'b000110;
 17'b00000010011001011 : data_comb = 6'b000101;
 17'b00000010011001100 : data_comb = 6'b000101;
 17'b00000010011001101 : data_comb = 6'b000101;
 17'b00000010011001110 : data_comb = 6'b000101;
 17'b00000010011001111 : data_comb = 6'b000101;
 17'b00000010011010000 : data_comb = 6'b000101;
 17'b00000010011010001 : data_comb = 6'b000101;
 17'b00000010011010010 : data_comb = 6'b000101;
 17'b00000010011010011 : data_comb = 6'b000101;
 17'b00000010011010100 : data_comb = 6'b000101;
 17'b00000010011010101 : data_comb = 6'b000101;
 17'b00000010011010110 : data_comb = 6'b000101;
 17'b00000010011010111 : data_comb = 6'b000101;
 17'b00000010011011000 : data_comb = 6'b000101;
 17'b00000010011011001 : data_comb = 6'b000101;
 17'b00000010011011010 : data_comb = 6'b000101;
 17'b00000010011011011 : data_comb = 6'b000101;
 17'b00000010011011100 : data_comb = 6'b000101;
 17'b00000010011011101 : data_comb = 6'b000101;
 17'b00000010011011110 : data_comb = 6'b000101;
 17'b00000010011011111 : data_comb = 6'b000101;
 17'b00000010011100000 : data_comb = 6'b000101;
 17'b00000010011100001 : data_comb = 6'b000101;
 17'b00000010011100010 : data_comb = 6'b111000;
 17'b00000010011100011 : data_comb = 6'b111000;
 17'b00000010011100100 : data_comb = 6'b111000;
 17'b00000010011100101 : data_comb = 6'b111000;
 17'b00000010011100110 : data_comb = 6'b111000;
 17'b00000010011100111 : data_comb = 6'b111000;
 17'b00000010011101000 : data_comb = 6'b111000;
 17'b00000010011101001 : data_comb = 6'b111000;
 17'b00000010011101010 : data_comb = 6'b111000;
 17'b00000010011101011 : data_comb = 6'b101000;
 17'b00000010011101100 : data_comb = 6'b101000;
 17'b00000010011101101 : data_comb = 6'b101000;
 17'b00000010011101110 : data_comb = 6'b000101;
 17'b00000010011101111 : data_comb = 6'b000101;
 17'b00000010011110000 : data_comb = 6'b000101;
 17'b00000010011110001 : data_comb = 6'b000101;
 17'b00000010011110010 : data_comb = 6'b000101;
 17'b00000010011110011 : data_comb = 6'b000101;
 17'b00000010011110100 : data_comb = 6'b000101;
 17'b00000010011110101 : data_comb = 6'b000101;
 17'b00000010011110110 : data_comb = 6'b000101;
 17'b00000010011110111 : data_comb = 6'b000101;
 17'b00000010011111000 : data_comb = 6'b000101;
 17'b00000010011111001 : data_comb = 6'b000101;
 17'b00000010011111010 : data_comb = 6'b101000;
 17'b00000010011111011 : data_comb = 6'b111000;
 17'b00000010011111100 : data_comb = 6'b111000;
 17'b00000010011111101 : data_comb = 6'b010101;
 17'b00000010011111110 : data_comb = 6'b000101;
 17'b00000010011111111 : data_comb = 6'b000101;
 17'b00000010100000000 : data_comb = 6'b111000;
 17'b00000010100000001 : data_comb = 6'b111000;
 17'b00000010100000010 : data_comb = 6'b111000;
 17'b00000010100000011 : data_comb = 6'b111000;
 17'b00000010100000100 : data_comb = 6'b111000;
 17'b00000010100000101 : data_comb = 6'b111000;
 17'b00000010100000110 : data_comb = 6'b111000;
 17'b00000010100000111 : data_comb = 6'b111000;
 17'b00000010100001000 : data_comb = 6'b111000;
 17'b00000010100001001 : data_comb = 6'b111000;
 17'b00000010100001010 : data_comb = 6'b111000;
 17'b00000010100001011 : data_comb = 6'b111000;
 17'b00000010100001100 : data_comb = 6'b111000;
 17'b00000010100001101 : data_comb = 6'b111000;
 17'b00000010100001110 : data_comb = 6'b101000;
 17'b00000010100001111 : data_comb = 6'b000101;
 17'b00000010100010000 : data_comb = 6'b000101;
 17'b00000010100010001 : data_comb = 6'b000101;
 17'b00000010100010010 : data_comb = 6'b000101;
 17'b00000010100010011 : data_comb = 6'b000101;
 17'b00000010100010100 : data_comb = 6'b000101;
 17'b00000010100010101 : data_comb = 6'b000101;
 17'b00000010100010110 : data_comb = 6'b000110;
 17'b00000010100010111 : data_comb = 6'b001010;
 17'b00000010100011000 : data_comb = 6'b001010;
 17'b00000010100011001 : data_comb = 6'b001010;
 17'b00000010100011010 : data_comb = 6'b001010;
 17'b00000010100011011 : data_comb = 6'b000110;
 17'b00000010100011100 : data_comb = 6'b000110;
 17'b00000010100011101 : data_comb = 6'b000110;
 17'b00000010100011110 : data_comb = 6'b000110;
 17'b00000010100011111 : data_comb = 6'b000101;
 17'b00000010100100000 : data_comb = 6'b000101;
 17'b00000010100100001 : data_comb = 6'b000101;
 17'b00000010100100010 : data_comb = 6'b000101;
 17'b00000010100100011 : data_comb = 6'b000101;
 17'b00000010100100100 : data_comb = 6'b000101;
 17'b00000010100100101 : data_comb = 6'b000101;
 17'b00000010100100110 : data_comb = 6'b000101;
 17'b00000010100100111 : data_comb = 6'b000101;
 17'b00000010100101000 : data_comb = 6'b000101;
 17'b00000010100101001 : data_comb = 6'b000101;
 17'b00000010100101010 : data_comb = 6'b000101;
 17'b00000010100101011 : data_comb = 6'b000101;
 17'b00000010100101100 : data_comb = 6'b000101;
 17'b00000010100101101 : data_comb = 6'b000101;
 17'b00000010100101110 : data_comb = 6'b000101;
 17'b00000010100101111 : data_comb = 6'b010101;
 17'b00000010100110000 : data_comb = 6'b010101;
 17'b00000010100110001 : data_comb = 6'b010101;
 17'b00000010100110010 : data_comb = 6'b111000;
 17'b00000010100110011 : data_comb = 6'b111000;
 17'b00000010100110100 : data_comb = 6'b111000;
 17'b00000010100110101 : data_comb = 6'b111000;
 17'b00000010100110110 : data_comb = 6'b111000;
 17'b00000010100110111 : data_comb = 6'b111000;
 17'b00000010100111000 : data_comb = 6'b111000;
 17'b00000010100111001 : data_comb = 6'b111000;
 17'b00000010100111010 : data_comb = 6'b111000;
 17'b00000010100111011 : data_comb = 6'b000101;
 17'b00000010100111100 : data_comb = 6'b000101;
 17'b00000010100111101 : data_comb = 6'b000101;
 17'b00000010100111110 : data_comb = 6'b000101;
 17'b00000010100111111 : data_comb = 6'b000101;
 17'b00000010101000000 : data_comb = 6'b000101;
 17'b00000010101000001 : data_comb = 6'b000101;
 17'b00000010101000010 : data_comb = 6'b000101;
 17'b00000010101000011 : data_comb = 6'b000101;
 17'b00000010101000100 : data_comb = 6'b000101;
 17'b00000010101000101 : data_comb = 6'b000101;
 17'b00000010101000110 : data_comb = 6'b000101;
 17'b00000010101000111 : data_comb = 6'b000101;
 17'b00000010101001000 : data_comb = 6'b000101;
 17'b00000010101001001 : data_comb = 6'b000101;
 17'b00000010101001010 : data_comb = 6'b111000;
 17'b00000010101001011 : data_comb = 6'b111000;
 17'b00000010101001100 : data_comb = 6'b111000;
 17'b00000010101001101 : data_comb = 6'b111000;
 17'b00000010101001110 : data_comb = 6'b000101;
 17'b00000010101001111 : data_comb = 6'b000101;
 17'b00000010101010000 : data_comb = 6'b000101;
 17'b00000010101010001 : data_comb = 6'b000101;
 17'b00000010101010010 : data_comb = 6'b000101;
 17'b00000010101010011 : data_comb = 6'b010101;
 17'b00000010101010100 : data_comb = 6'b111000;
 17'b00000010101010101 : data_comb = 6'b111000;
 17'b00000010101010110 : data_comb = 6'b111000;
 17'b00000010101010111 : data_comb = 6'b111000;
 17'b00000010101011000 : data_comb = 6'b111000;
 17'b00000010101011001 : data_comb = 6'b111000;
 17'b00000010101011010 : data_comb = 6'b111000;
 17'b00000010101011011 : data_comb = 6'b111000;
 17'b00000010101011100 : data_comb = 6'b111000;
 17'b00000010101011101 : data_comb = 6'b111000;
 17'b00000010101011110 : data_comb = 6'b111000;
 17'b00000010101011111 : data_comb = 6'b111000;
 17'b00000010101100000 : data_comb = 6'b111000;
 17'b00000010101100001 : data_comb = 6'b000101;
 17'b00000010101100010 : data_comb = 6'b000101;
 17'b00000010101100011 : data_comb = 6'b000101;
 17'b00000010101100100 : data_comb = 6'b000101;
 17'b00000010101100101 : data_comb = 6'b000101;
 17'b00000010101100110 : data_comb = 6'b000101;
 17'b00000010101100111 : data_comb = 6'b000101;
 17'b00000010101101000 : data_comb = 6'b000110;
 17'b00000010101101001 : data_comb = 6'b001010;
 17'b00000010101101010 : data_comb = 6'b001010;
 17'b00000010101101011 : data_comb = 6'b001010;
 17'b00000010101101100 : data_comb = 6'b001010;
 17'b00000010101101101 : data_comb = 6'b001010;
 17'b00000010101101110 : data_comb = 6'b000110;
 17'b00000010101101111 : data_comb = 6'b000101;
 17'b00000010101110000 : data_comb = 6'b000101;
 17'b00000010101110001 : data_comb = 6'b000101;
 17'b00000010101110010 : data_comb = 6'b000101;
 17'b00000010101110011 : data_comb = 6'b000101;
 17'b00000010101110100 : data_comb = 6'b000101;
 17'b00000010101110101 : data_comb = 6'b000101;
 17'b00000010101110110 : data_comb = 6'b000101;
 17'b00000010101110111 : data_comb = 6'b000101;
 17'b00000010101111000 : data_comb = 6'b000101;
 17'b00000010101111001 : data_comb = 6'b000101;
 17'b00000010101111010 : data_comb = 6'b000101;
 17'b00000010101111011 : data_comb = 6'b000101;
 17'b00000010101111100 : data_comb = 6'b000101;
 17'b00000010101111101 : data_comb = 6'b101000;
 17'b00000010101111110 : data_comb = 6'b101000;
 17'b00000010101111111 : data_comb = 6'b111000;
 17'b00000010110000000 : data_comb = 6'b111000;
 17'b00000010110000001 : data_comb = 6'b111000;
 17'b00000010110000010 : data_comb = 6'b111000;
 17'b00000010110000011 : data_comb = 6'b111000;
 17'b00000010110000100 : data_comb = 6'b111000;
 17'b00000010110000101 : data_comb = 6'b111000;
 17'b00000010110000110 : data_comb = 6'b010101;
 17'b00000010110000111 : data_comb = 6'b010101;
 17'b00000010110001000 : data_comb = 6'b100101;
 17'b00000010110001001 : data_comb = 6'b111000;
 17'b00000010110001010 : data_comb = 6'b111000;
 17'b00000010110001011 : data_comb = 6'b101000;
 17'b00000010110001100 : data_comb = 6'b010101;
 17'b00000010110001101 : data_comb = 6'b000101;
 17'b00000010110001110 : data_comb = 6'b000101;
 17'b00000010110001111 : data_comb = 6'b000101;
 17'b00000010110010000 : data_comb = 6'b000101;
 17'b00000010110010001 : data_comb = 6'b000101;
 17'b00000010110010010 : data_comb = 6'b000101;
 17'b00000010110010011 : data_comb = 6'b000101;
 17'b00000010110010100 : data_comb = 6'b000101;
 17'b00000010110010101 : data_comb = 6'b000101;
 17'b00000010110010110 : data_comb = 6'b000101;
 17'b00000010110010111 : data_comb = 6'b000101;
 17'b00000010110011000 : data_comb = 6'b101000;
 17'b00000010110011001 : data_comb = 6'b101000;
 17'b00000010110011010 : data_comb = 6'b111000;
 17'b00000010110011011 : data_comb = 6'b111000;
 17'b00000010110011100 : data_comb = 6'b111000;
 17'b00000010110011101 : data_comb = 6'b111000;
 17'b00000010110011110 : data_comb = 6'b101000;
 17'b00000010110011111 : data_comb = 6'b101000;
 17'b00000010110100000 : data_comb = 6'b000101;
 17'b00000010110100001 : data_comb = 6'b000101;
 17'b00000010110100010 : data_comb = 6'b000101;
 17'b00000010110100011 : data_comb = 6'b111000;
 17'b00000010110100100 : data_comb = 6'b111000;
 17'b00000010110100101 : data_comb = 6'b111000;
 17'b00000010110100110 : data_comb = 6'b111000;
 17'b00000010110100111 : data_comb = 6'b111000;
 17'b00000010110101000 : data_comb = 6'b010101;
 17'b00000010110101001 : data_comb = 6'b010101;
 17'b00000010110101010 : data_comb = 6'b010101;
 17'b00000010110101011 : data_comb = 6'b010101;
 17'b00000010110101100 : data_comb = 6'b111000;
 17'b00000010110101101 : data_comb = 6'b111000;
 17'b00000010110101110 : data_comb = 6'b111000;
 17'b00000010110101111 : data_comb = 6'b111000;
 17'b00000010110110000 : data_comb = 6'b111000;
 17'b00000010110110001 : data_comb = 6'b101000;
 17'b00000010110110010 : data_comb = 6'b101001;
 17'b00000010110110011 : data_comb = 6'b101001;
 17'b00000010110110100 : data_comb = 6'b000101;
 17'b00000010110110101 : data_comb = 6'b000101;
 17'b00000010110110110 : data_comb = 6'b000101;
 17'b00000010110110111 : data_comb = 6'b000101;
 17'b00000010110111000 : data_comb = 6'b000101;
 17'b00000010110111001 : data_comb = 6'b000101;
 17'b00000010110111010 : data_comb = 6'b000101;
 17'b00000010110111011 : data_comb = 6'b000101;
 17'b00000010110111100 : data_comb = 6'b000101;
 17'b00000010110111101 : data_comb = 6'b000101;
 17'b00000010110111110 : data_comb = 6'b000101;
 17'b00000010110111111 : data_comb = 6'b000101;
 17'b00000010111000000 : data_comb = 6'b000101;
 17'b00000010111000001 : data_comb = 6'b000101;
 17'b00000010111000010 : data_comb = 6'b000101;
 17'b00000010111000011 : data_comb = 6'b000101;
 17'b00000010111000100 : data_comb = 6'b000101;
 17'b00000010111000101 : data_comb = 6'b000101;
 17'b00000010111000110 : data_comb = 6'b000101;
 17'b00000010111000111 : data_comb = 6'b000101;
 17'b00000010111001000 : data_comb = 6'b000101;
 17'b00000010111001001 : data_comb = 6'b000101;
 17'b00000010111001010 : data_comb = 6'b000101;
 17'b00000010111001011 : data_comb = 6'b000101;
 17'b00000010111001100 : data_comb = 6'b010101;
 17'b00000010111001101 : data_comb = 6'b111000;
 17'b00000010111001110 : data_comb = 6'b111000;
 17'b00000010111001111 : data_comb = 6'b111000;
 17'b00000010111010000 : data_comb = 6'b111000;
 17'b00000010111010001 : data_comb = 6'b111000;
 17'b00000010111010010 : data_comb = 6'b111000;
 17'b00000010111010011 : data_comb = 6'b111000;
 17'b00000010111010100 : data_comb = 6'b111000;
 17'b00000010111010101 : data_comb = 6'b101000;
 17'b00000010111010110 : data_comb = 6'b000101;
 17'b00000010111010111 : data_comb = 6'b000101;
 17'b00000010111011000 : data_comb = 6'b010101;
 17'b00000010111011001 : data_comb = 6'b111000;
 17'b00000010111011010 : data_comb = 6'b111000;
 17'b00000010111011011 : data_comb = 6'b111000;
 17'b00000010111011100 : data_comb = 6'b101000;
 17'b00000010111011101 : data_comb = 6'b000101;
 17'b00000010111011110 : data_comb = 6'b000101;
 17'b00000010111011111 : data_comb = 6'b000101;
 17'b00000010111100000 : data_comb = 6'b000101;
 17'b00000010111100001 : data_comb = 6'b101001;
 17'b00000010111100010 : data_comb = 6'b111000;
 17'b00000010111100011 : data_comb = 6'b111000;
 17'b00000010111100100 : data_comb = 6'b000101;
 17'b00000010111100101 : data_comb = 6'b000101;
 17'b00000010111100110 : data_comb = 6'b000101;
 17'b00000010111100111 : data_comb = 6'b101000;
 17'b00000010111101000 : data_comb = 6'b111000;
 17'b00000010111101001 : data_comb = 6'b111000;
 17'b00000010111101010 : data_comb = 6'b111000;
 17'b00000010111101011 : data_comb = 6'b111000;
 17'b00000010111101100 : data_comb = 6'b111000;
 17'b00000010111101101 : data_comb = 6'b111000;
 17'b00000010111101110 : data_comb = 6'b111000;
 17'b00000010111101111 : data_comb = 6'b111000;
 17'b00000010111110000 : data_comb = 6'b000101;
 17'b00000010111110001 : data_comb = 6'b000101;
 17'b00000010111110010 : data_comb = 6'b000101;
 17'b00000010111110011 : data_comb = 6'b000101;
 17'b00000010111110100 : data_comb = 6'b000101;
 17'b00000010111110101 : data_comb = 6'b000101;
 17'b00000010111110110 : data_comb = 6'b000101;
 17'b00000010111110111 : data_comb = 6'b000101;
 17'b00000010111111000 : data_comb = 6'b000101;
 17'b00000010111111001 : data_comb = 6'b000101;
 17'b00000010111111010 : data_comb = 6'b000101;
 17'b00000010111111011 : data_comb = 6'b000101;
 17'b00000010111111100 : data_comb = 6'b101000;
 17'b00000010111111101 : data_comb = 6'b101000;
 17'b00000010111111110 : data_comb = 6'b101000;
 17'b00000010111111111 : data_comb = 6'b101000;
 17'b00000011000000000 : data_comb = 6'b111000;
 17'b00000011000000001 : data_comb = 6'b111000;
 17'b00000011000000010 : data_comb = 6'b111000;
 17'b00000011000000011 : data_comb = 6'b111000;
 17'b00000011000000100 : data_comb = 6'b010101;
 17'b00000011000000101 : data_comb = 6'b000101;
 17'b00000011000000110 : data_comb = 6'b000101;
 17'b00000011000000111 : data_comb = 6'b000101;
 17'b00000011000001000 : data_comb = 6'b000101;
 17'b00000011000001001 : data_comb = 6'b000101;
 17'b00000011000001010 : data_comb = 6'b000101;
 17'b00000011000001011 : data_comb = 6'b000101;
 17'b00000011000001100 : data_comb = 6'b000101;
 17'b00000011000001101 : data_comb = 6'b000101;
 17'b00000011000001110 : data_comb = 6'b000101;
 17'b00000011000001111 : data_comb = 6'b000101;
 17'b00000011000010000 : data_comb = 6'b000101;
 17'b00000011000010001 : data_comb = 6'b000101;
 17'b00000011000010010 : data_comb = 6'b000101;
 17'b00000011000010011 : data_comb = 6'b000101;
 17'b00000011000010100 : data_comb = 6'b000101;
 17'b00000011000010101 : data_comb = 6'b000101;
 17'b00000011000010110 : data_comb = 6'b000101;
 17'b00000011000010111 : data_comb = 6'b000101;
 17'b00000011000011000 : data_comb = 6'b000101;
 17'b00000011000011001 : data_comb = 6'b000101;
 17'b00000011000011010 : data_comb = 6'b000101;
 17'b00000011000011011 : data_comb = 6'b000101;
 17'b00000011000011100 : data_comb = 6'b000101;
 17'b00000011000011101 : data_comb = 6'b000101;
 17'b00000011000011110 : data_comb = 6'b000110;
 17'b00000011000011111 : data_comb = 6'b000101;
 17'b00000011000100000 : data_comb = 6'b000101;
 17'b00000011000100001 : data_comb = 6'b000101;
 17'b00000011000100010 : data_comb = 6'b000101;
 17'b00000011000100011 : data_comb = 6'b000110;
 17'b00000011000100100 : data_comb = 6'b000101;
 17'b00000011000100101 : data_comb = 6'b000101;
 17'b00000011000100110 : data_comb = 6'b000101;
 17'b00000011000100111 : data_comb = 6'b000101;
 17'b00000011000101000 : data_comb = 6'b000101;
 17'b00000011000101001 : data_comb = 6'b000101;
 17'b00000011000101010 : data_comb = 6'b000101;
 17'b00000011000101011 : data_comb = 6'b000101;
 17'b00000011000101100 : data_comb = 6'b000101;
 17'b00000011000101101 : data_comb = 6'b000101;
 17'b00000011000101110 : data_comb = 6'b000101;
 17'b00000011000101111 : data_comb = 6'b000101;
 17'b00000011000110000 : data_comb = 6'b101001;
 17'b00000011000110001 : data_comb = 6'b111000;
 17'b00000011000110010 : data_comb = 6'b111000;
 17'b00000011000110011 : data_comb = 6'b111000;
 17'b00000011000110100 : data_comb = 6'b111000;
 17'b00000011000110101 : data_comb = 6'b010101;
 17'b00000011000110110 : data_comb = 6'b000101;
 17'b00000011000110111 : data_comb = 6'b000101;
 17'b00000011000111000 : data_comb = 6'b000101;
 17'b00000011000111001 : data_comb = 6'b000101;
 17'b00000011000111010 : data_comb = 6'b000101;
 17'b00000011000111011 : data_comb = 6'b111000;
 17'b00000011000111100 : data_comb = 6'b111000;
 17'b00000011000111101 : data_comb = 6'b111000;
 17'b00000011000111110 : data_comb = 6'b010101;
 17'b00000011000111111 : data_comb = 6'b000101;
 17'b00000011001000000 : data_comb = 6'b000101;
 17'b00000011001000001 : data_comb = 6'b000101;
 17'b00000011001000010 : data_comb = 6'b000101;
 17'b00000011001000011 : data_comb = 6'b000101;
 17'b00000011001000100 : data_comb = 6'b000101;
 17'b00000011001000101 : data_comb = 6'b000101;
 17'b00000011001000110 : data_comb = 6'b000101;
 17'b00000011001000111 : data_comb = 6'b000101;
 17'b00000011001001000 : data_comb = 6'b000101;
 17'b00000011001001001 : data_comb = 6'b000101;
 17'b00000011001001010 : data_comb = 6'b000101;
 17'b00000011001001011 : data_comb = 6'b000101;
 17'b00000011001001100 : data_comb = 6'b000101;
 17'b00000011001001101 : data_comb = 6'b000101;
 17'b00000011001001110 : data_comb = 6'b000101;
 17'b00000011001001111 : data_comb = 6'b000101;
 17'b00000011001010000 : data_comb = 6'b010101;
 17'b00000011001010001 : data_comb = 6'b010101;
 17'b00000011001010010 : data_comb = 6'b010101;
 17'b00000011001010011 : data_comb = 6'b010101;
 17'b00000011001010100 : data_comb = 6'b000101;
 17'b00000011001010101 : data_comb = 6'b000101;
 17'b00000011001010110 : data_comb = 6'b000101;
 17'b00000011001010111 : data_comb = 6'b000101;
 17'b00000011001011000 : data_comb = 6'b000101;
 17'b00000011001011001 : data_comb = 6'b000101;
 17'b00000011001011010 : data_comb = 6'b000101;
 17'b00000011001011011 : data_comb = 6'b000101;
 17'b00000011001011100 : data_comb = 6'b000101;
 17'b00000011001011101 : data_comb = 6'b000101;
 17'b00000011001011110 : data_comb = 6'b000101;
 17'b00000011001011111 : data_comb = 6'b000101;
 17'b00000011001100000 : data_comb = 6'b000101;
 17'b00000011001100001 : data_comb = 6'b101000;
 17'b00000011001100010 : data_comb = 6'b101000;
 17'b00000011001100011 : data_comb = 6'b000101;
 17'b00000011001100100 : data_comb = 6'b000101;
 17'b00000011001100101 : data_comb = 6'b000101;
 17'b00000011001100110 : data_comb = 6'b000101;
 17'b00000011001100111 : data_comb = 6'b000101;
 17'b00000011001101000 : data_comb = 6'b000101;
 17'b00000011001101001 : data_comb = 6'b000101;
 17'b00000011001101010 : data_comb = 6'b000101;
 17'b00000011001101011 : data_comb = 6'b000101;
 17'b00000011001101100 : data_comb = 6'b000101;
 17'b00000011001101101 : data_comb = 6'b000101;
 17'b00000011001101110 : data_comb = 6'b000101;
 17'b00000011001101111 : data_comb = 6'b000101;
 17'b00000011001110000 : data_comb = 6'b000101;
 17'b00000011001110001 : data_comb = 6'b000101;
 17'b00000011001110010 : data_comb = 6'b000101;
 17'b00000011001110011 : data_comb = 6'b000101;
 17'b00000011001110100 : data_comb = 6'b000101;
 17'b00000011001110101 : data_comb = 6'b000101;
 17'b00000011001110110 : data_comb = 6'b000101;
 17'b00000011001110111 : data_comb = 6'b000101;
 17'b00000011001111000 : data_comb = 6'b000101;
 17'b00000011001111001 : data_comb = 6'b000101;
 17'b00000011001111010 : data_comb = 6'b000101;
 17'b00000011001111011 : data_comb = 6'b000101;
 17'b00000011001111100 : data_comb = 6'b000101;
 17'b00000011001111101 : data_comb = 6'b000101;
 17'b00000011001111110 : data_comb = 6'b000101;
 17'b00000011001111111 : data_comb = 6'b000101;
 17'b00000011010000000 : data_comb = 6'b101000;
 17'b00000011010000001 : data_comb = 6'b111000;
 17'b00000011010000010 : data_comb = 6'b111000;
 17'b00000011010000011 : data_comb = 6'b111000;
 17'b00000011010000100 : data_comb = 6'b111000;
 17'b00000011010000101 : data_comb = 6'b111000;
 17'b00000011010000110 : data_comb = 6'b000101;
 17'b00000011010000111 : data_comb = 6'b000101;
 17'b00000011010001000 : data_comb = 6'b000101;
 17'b00000011010001001 : data_comb = 6'b000101;
 17'b00000011010001010 : data_comb = 6'b000101;
 17'b00000011010001011 : data_comb = 6'b000101;
 17'b00000011010001100 : data_comb = 6'b000101;
 17'b00000011010001101 : data_comb = 6'b000101;
 17'b00000011010001110 : data_comb = 6'b000101;
 17'b00000011010001111 : data_comb = 6'b000101;
 17'b00000011010010000 : data_comb = 6'b000101;
 17'b00000011010010001 : data_comb = 6'b000101;
 17'b00000011010010010 : data_comb = 6'b000101;
 17'b00000011010010011 : data_comb = 6'b000101;
 17'b00000011010010100 : data_comb = 6'b000101;
 17'b00000011010010101 : data_comb = 6'b000101;
 17'b00000011010010110 : data_comb = 6'b000101;
 17'b00000011010010111 : data_comb = 6'b000101;
 17'b00000011010011000 : data_comb = 6'b000101;
 17'b00000011010011001 : data_comb = 6'b000101;
 17'b00000011010011010 : data_comb = 6'b000101;
 17'b00000011010011011 : data_comb = 6'b000101;
 17'b00000011010011100 : data_comb = 6'b000101;
 17'b00000011010011101 : data_comb = 6'b000101;
 17'b00000011010011110 : data_comb = 6'b000101;
 17'b00000011010011111 : data_comb = 6'b000101;
 17'b00000011010100000 : data_comb = 6'b000101;
 17'b00000011010100001 : data_comb = 6'b000101;
 17'b00000011010100010 : data_comb = 6'b000101;
 17'b00000011010100011 : data_comb = 6'b000101;
 17'b00000011010100100 : data_comb = 6'b000101;
 17'b00000011010100101 : data_comb = 6'b000101;
 17'b00000011010100110 : data_comb = 6'b000101;
 17'b00000011010100111 : data_comb = 6'b000101;
 17'b00000011010101000 : data_comb = 6'b000101;
 17'b00000011010101001 : data_comb = 6'b000101;
 17'b00000011010101010 : data_comb = 6'b000101;
 17'b00000011010101011 : data_comb = 6'b000101;
 17'b00000011010101100 : data_comb = 6'b000101;
 17'b00000011010101101 : data_comb = 6'b000101;
 17'b00000011010101110 : data_comb = 6'b000101;
 17'b00000011010101111 : data_comb = 6'b000101;
 17'b00000011010110000 : data_comb = 6'b111000;
 17'b00000011010110001 : data_comb = 6'b111000;
 17'b00000011010110010 : data_comb = 6'b111000;
 17'b00000011010110011 : data_comb = 6'b111000;
 17'b00000011010110100 : data_comb = 6'b010101;
 17'b00000011010110101 : data_comb = 6'b000101;
 17'b00000011010110110 : data_comb = 6'b000101;
 17'b00000011010110111 : data_comb = 6'b000101;
 17'b00000011010111000 : data_comb = 6'b000101;
 17'b00000011010111001 : data_comb = 6'b000101;
 17'b00000011010111010 : data_comb = 6'b000101;
 17'b00000011010111011 : data_comb = 6'b000101;
 17'b00000011010111100 : data_comb = 6'b000101;
 17'b00000011010111101 : data_comb = 6'b000101;
 17'b00000011010111110 : data_comb = 6'b000101;
 17'b00000011010111111 : data_comb = 6'b000101;
 17'b00000011011000000 : data_comb = 6'b000101;
 17'b00000011011000001 : data_comb = 6'b000101;
 17'b00000011011000010 : data_comb = 6'b000101;
 17'b00000011011000011 : data_comb = 6'b000101;
 17'b00000011011000100 : data_comb = 6'b000101;
 17'b00000011011000101 : data_comb = 6'b000101;
 17'b00000011011000110 : data_comb = 6'b000101;
 17'b00000011011000111 : data_comb = 6'b000101;
 17'b00000011011001000 : data_comb = 6'b000101;
 17'b00000011011001001 : data_comb = 6'b000101;
 17'b00000011011001010 : data_comb = 6'b000101;
 17'b00000011011001011 : data_comb = 6'b000101;
 17'b00000011011001100 : data_comb = 6'b000101;
 17'b00000011011001101 : data_comb = 6'b000101;
 17'b00000011011001110 : data_comb = 6'b000101;
 17'b00000011011001111 : data_comb = 6'b010101;
 17'b00000011011010000 : data_comb = 6'b111000;
 17'b00000011011010001 : data_comb = 6'b111000;
 17'b00000011011010010 : data_comb = 6'b111000;
 17'b00000011011010011 : data_comb = 6'b111000;
 17'b00000011011010100 : data_comb = 6'b111000;
 17'b00000011011010101 : data_comb = 6'b111000;
 17'b00000011011010110 : data_comb = 6'b010101;
 17'b00000011011010111 : data_comb = 6'b000101;
 17'b00000011011011000 : data_comb = 6'b000101;
 17'b00000011011011001 : data_comb = 6'b000101;
 17'b00000011011011010 : data_comb = 6'b000101;
 17'b00000011011011011 : data_comb = 6'b000101;
 17'b00000011011011100 : data_comb = 6'b000101;
 17'b00000011011011101 : data_comb = 6'b000101;
 17'b00000011011011110 : data_comb = 6'b000101;
 17'b00000011011011111 : data_comb = 6'b000101;
 17'b00000011011100000 : data_comb = 6'b000101;
 17'b00000011011100001 : data_comb = 6'b000101;
 17'b00000011011100010 : data_comb = 6'b000101;
 17'b00000011011100011 : data_comb = 6'b000101;
 17'b00000011011100100 : data_comb = 6'b000101;
 17'b00000011011100101 : data_comb = 6'b000101;
 17'b00000011011100110 : data_comb = 6'b000101;
 17'b00000011011100111 : data_comb = 6'b000101;
 17'b00000011011101000 : data_comb = 6'b000101;
 17'b00000011011101001 : data_comb = 6'b101001;
 17'b00000011011101010 : data_comb = 6'b011001;
 17'b00000011011101011 : data_comb = 6'b000101;
 17'b00000011011101100 : data_comb = 6'b000101;
 17'b00000011011101101 : data_comb = 6'b000101;
 17'b00000011011101110 : data_comb = 6'b000101;
 17'b00000011011101111 : data_comb = 6'b000101;
 17'b00000011011110000 : data_comb = 6'b000101;
 17'b00000011011110001 : data_comb = 6'b000101;
 17'b00000011011110010 : data_comb = 6'b000101;
 17'b00000011011110011 : data_comb = 6'b000101;
 17'b00000011011110100 : data_comb = 6'b000101;
 17'b00000011011110101 : data_comb = 6'b000101;
 17'b00000011011110110 : data_comb = 6'b000101;
 17'b00000011011110111 : data_comb = 6'b000101;
 17'b00000011011111000 : data_comb = 6'b000101;
 17'b00000011011111001 : data_comb = 6'b000101;
 17'b00000011011111010 : data_comb = 6'b000101;
 17'b00000011011111011 : data_comb = 6'b000101;
 17'b00000011011111100 : data_comb = 6'b000101;
 17'b00000011011111101 : data_comb = 6'b010101;
 17'b00000011011111110 : data_comb = 6'b111000;
 17'b00000011011111111 : data_comb = 6'b111000;
 17'b00000011100000000 : data_comb = 6'b111000;
 17'b00000011100000001 : data_comb = 6'b111000;
 17'b00000011100000010 : data_comb = 6'b111000;
 17'b00000011100000011 : data_comb = 6'b111000;
 17'b00000011100000100 : data_comb = 6'b111000;
 17'b00000011100000101 : data_comb = 6'b101000;
 17'b00000011100000110 : data_comb = 6'b010101;
 17'b00000011100000111 : data_comb = 6'b000101;
 17'b00000011100001000 : data_comb = 6'b000101;
 17'b00000011100001001 : data_comb = 6'b000101;
 17'b00000011100001010 : data_comb = 6'b000101;
 17'b00000011100001011 : data_comb = 6'b000101;
 17'b00000011100001100 : data_comb = 6'b000101;
 17'b00000011100001101 : data_comb = 6'b000101;
 17'b00000011100001110 : data_comb = 6'b000101;
 17'b00000011100001111 : data_comb = 6'b000101;
 17'b00000011100010000 : data_comb = 6'b000101;
 17'b00000011100010001 : data_comb = 6'b000101;
 17'b00000011100010010 : data_comb = 6'b000101;
 17'b00000011100010011 : data_comb = 6'b000101;
 17'b00000011100010100 : data_comb = 6'b000101;
 17'b00000011100010101 : data_comb = 6'b000101;
 17'b00000011100010110 : data_comb = 6'b000101;
 17'b00000011100010111 : data_comb = 6'b000101;
 17'b00000011100011000 : data_comb = 6'b000101;
 17'b00000011100011001 : data_comb = 6'b000101;
 17'b00000011100011010 : data_comb = 6'b000101;
 17'b00000011100011011 : data_comb = 6'b000101;
 17'b00000011100011100 : data_comb = 6'b000101;
 17'b00000011100011101 : data_comb = 6'b000101;
 17'b00000011100011110 : data_comb = 6'b000101;
 17'b00000011100011111 : data_comb = 6'b000101;
 17'b00000011100100000 : data_comb = 6'b101000;
 17'b00000011100100001 : data_comb = 6'b111000;
 17'b00000011100100010 : data_comb = 6'b111000;
 17'b00000011100100011 : data_comb = 6'b111000;
 17'b00000011100100100 : data_comb = 6'b111000;
 17'b00000011100100101 : data_comb = 6'b111000;
 17'b00000011100100110 : data_comb = 6'b111000;
 17'b00000011100100111 : data_comb = 6'b010101;
 17'b00000011100101000 : data_comb = 6'b000101;
 17'b00000011100101001 : data_comb = 6'b010101;
 17'b00000011100101010 : data_comb = 6'b010101;
 17'b00000011100101011 : data_comb = 6'b000101;
 17'b00000011100101100 : data_comb = 6'b000101;
 17'b00000011100101101 : data_comb = 6'b000101;
 17'b00000011100101110 : data_comb = 6'b000101;
 17'b00000011100101111 : data_comb = 6'b000101;
 17'b00000011100110000 : data_comb = 6'b000101;
 17'b00000011100110001 : data_comb = 6'b000101;
 17'b00000011100110010 : data_comb = 6'b000101;
 17'b00000011100110011 : data_comb = 6'b000101;
 17'b00000011100110100 : data_comb = 6'b000101;
 17'b00000011100110101 : data_comb = 6'b000101;
 17'b00000011100110110 : data_comb = 6'b000101;
 17'b00000011100110111 : data_comb = 6'b000101;
 17'b00000011100111000 : data_comb = 6'b111000;
 17'b00000011100111001 : data_comb = 6'b111000;
 17'b00000011100111010 : data_comb = 6'b111000;
 17'b00000011100111011 : data_comb = 6'b101000;
 17'b00000011100111100 : data_comb = 6'b000101;
 17'b00000011100111101 : data_comb = 6'b000101;
 17'b00000011100111110 : data_comb = 6'b000101;
 17'b00000011100111111 : data_comb = 6'b000101;
 17'b00000011101000000 : data_comb = 6'b000101;
 17'b00000011101000001 : data_comb = 6'b000101;
 17'b00000011101000010 : data_comb = 6'b000101;
 17'b00000011101000011 : data_comb = 6'b000101;
 17'b00000011101000100 : data_comb = 6'b000101;
 17'b00000011101000101 : data_comb = 6'b000101;
 17'b00000011101000110 : data_comb = 6'b000101;
 17'b00000011101000111 : data_comb = 6'b000101;
 17'b00000011101001000 : data_comb = 6'b000101;
 17'b00000011101001001 : data_comb = 6'b000101;
 17'b00000011101001010 : data_comb = 6'b000101;
 17'b00000011101001011 : data_comb = 6'b000101;
 17'b00000011101001100 : data_comb = 6'b000101;
 17'b00000011101001101 : data_comb = 6'b000101;
 17'b00000011101001110 : data_comb = 6'b010101;
 17'b00000011101001111 : data_comb = 6'b010101;
 17'b00000011101010000 : data_comb = 6'b111000;
 17'b00000011101010001 : data_comb = 6'b111000;
 17'b00000011101010010 : data_comb = 6'b111000;
 17'b00000011101010011 : data_comb = 6'b111000;
 17'b00000011101010100 : data_comb = 6'b101000;
 17'b00000011101010101 : data_comb = 6'b010101;
 17'b00000011101010110 : data_comb = 6'b000101;
 17'b00000011101010111 : data_comb = 6'b000101;
 17'b00000011101011000 : data_comb = 6'b000101;
 17'b00000011101011001 : data_comb = 6'b000101;
 17'b00000011101011010 : data_comb = 6'b000101;
 17'b00000011101011011 : data_comb = 6'b000101;
 17'b00000011101011100 : data_comb = 6'b000101;
 17'b00000011101011101 : data_comb = 6'b000101;
 17'b00000011101011110 : data_comb = 6'b000101;
 17'b00000011101011111 : data_comb = 6'b000101;
 17'b00000011101100000 : data_comb = 6'b000101;
 17'b00000011101100001 : data_comb = 6'b000101;
 17'b00000011101100010 : data_comb = 6'b000101;
 17'b00000011101100011 : data_comb = 6'b000101;
 17'b00000011101100100 : data_comb = 6'b000101;
 17'b00000011101100101 : data_comb = 6'b000101;
 17'b00000011101100110 : data_comb = 6'b000101;
 17'b00000011101100111 : data_comb = 6'b000101;
 17'b00000011101101000 : data_comb = 6'b000101;
 17'b00000011101101001 : data_comb = 6'b000101;
 17'b00000011101101010 : data_comb = 6'b000101;
 17'b00000011101101011 : data_comb = 6'b000101;
 17'b00000011101101100 : data_comb = 6'b000101;
 17'b00000011101101101 : data_comb = 6'b000101;
 17'b00000011101101110 : data_comb = 6'b000101;
 17'b00000011101101111 : data_comb = 6'b000101;
 17'b00000011101110000 : data_comb = 6'b010101;
 17'b00000011101110001 : data_comb = 6'b111000;
 17'b00000011101110010 : data_comb = 6'b111000;
 17'b00000011101110011 : data_comb = 6'b111000;
 17'b00000011101110100 : data_comb = 6'b111000;
 17'b00000011101110101 : data_comb = 6'b111000;
 17'b00000011101110110 : data_comb = 6'b111000;
 17'b00000011101110111 : data_comb = 6'b111000;
 17'b00000011101111000 : data_comb = 6'b101000;
 17'b00000011101111001 : data_comb = 6'b111000;
 17'b00000011101111010 : data_comb = 6'b111000;
 17'b00000011101111011 : data_comb = 6'b101000;
 17'b00000011101111100 : data_comb = 6'b000101;
 17'b00000011101111101 : data_comb = 6'b000101;
 17'b00000011101111110 : data_comb = 6'b000101;
 17'b00000011101111111 : data_comb = 6'b000101;
 17'b00000011110000000 : data_comb = 6'b000101;
 17'b00000011110000001 : data_comb = 6'b000101;
 17'b00000011110000010 : data_comb = 6'b000101;
 17'b00000011110000011 : data_comb = 6'b000101;
 17'b00000011110000100 : data_comb = 6'b000101;
 17'b00000011110000101 : data_comb = 6'b000101;
 17'b00000011110000110 : data_comb = 6'b000101;
 17'b00000011110000111 : data_comb = 6'b101000;
 17'b00000011110001000 : data_comb = 6'b111000;
 17'b00000011110001001 : data_comb = 6'b111000;
 17'b00000011110001010 : data_comb = 6'b111000;
 17'b00000011110001011 : data_comb = 6'b101000;
 17'b00000011110001100 : data_comb = 6'b000101;
 17'b00000011110001101 : data_comb = 6'b000101;
 17'b00000011110001110 : data_comb = 6'b000101;
 17'b00000011110001111 : data_comb = 6'b000101;
 17'b00000011110010000 : data_comb = 6'b000101;
 17'b00000011110010001 : data_comb = 6'b000101;
 17'b00000011110010010 : data_comb = 6'b000101;
 17'b00000011110010011 : data_comb = 6'b000101;
 17'b00000011110010100 : data_comb = 6'b000101;
 17'b00000011110010101 : data_comb = 6'b000101;
 17'b00000011110010110 : data_comb = 6'b000101;
 17'b00000011110010111 : data_comb = 6'b000101;
 17'b00000011110011000 : data_comb = 6'b000101;
 17'b00000011110011001 : data_comb = 6'b000101;
 17'b00000011110011010 : data_comb = 6'b000101;
 17'b00000011110011011 : data_comb = 6'b000101;
 17'b00000011110011100 : data_comb = 6'b000101;
 17'b00000011110011101 : data_comb = 6'b000101;
 17'b00000011110011110 : data_comb = 6'b000101;
 17'b00000011110011111 : data_comb = 6'b000101;
 17'b00000011110100000 : data_comb = 6'b000101;
 17'b00000011110100001 : data_comb = 6'b000101;
 17'b00000011110100010 : data_comb = 6'b000101;
 17'b00000011110100011 : data_comb = 6'b000101;
 17'b00000011110100100 : data_comb = 6'b000101;
 17'b00000011110100101 : data_comb = 6'b000101;
 17'b00000011110100110 : data_comb = 6'b000101;
 17'b00000011110100111 : data_comb = 6'b000101;
 17'b00000011110101000 : data_comb = 6'b000101;
 17'b00000011110101001 : data_comb = 6'b000101;
 17'b00000011110101010 : data_comb = 6'b000101;
 17'b00000011110101011 : data_comb = 6'b000101;
 17'b00000011110101100 : data_comb = 6'b000101;
 17'b00000011110101101 : data_comb = 6'b000101;
 17'b00000011110101110 : data_comb = 6'b000101;
 17'b00000011110101111 : data_comb = 6'b000101;
 17'b00000011110110000 : data_comb = 6'b000101;
 17'b00000011110110001 : data_comb = 6'b000101;
 17'b00000011110110010 : data_comb = 6'b000101;
 17'b00000011110110011 : data_comb = 6'b000101;
 17'b00000011110110100 : data_comb = 6'b000101;
 17'b00000011110110101 : data_comb = 6'b000101;
 17'b00000011110110110 : data_comb = 6'b000101;
 17'b00000011110110111 : data_comb = 6'b000101;
 17'b00000011110111000 : data_comb = 6'b000101;
 17'b00000011110111001 : data_comb = 6'b000101;
 17'b00000011110111010 : data_comb = 6'b000101;
 17'b00000011110111011 : data_comb = 6'b000101;
 17'b00000011110111100 : data_comb = 6'b000101;
 17'b00000011110111101 : data_comb = 6'b000101;
 17'b00000011110111110 : data_comb = 6'b000101;
 17'b00000011110111111 : data_comb = 6'b000101;
 17'b00000011111000000 : data_comb = 6'b000101;
 17'b00000011111000001 : data_comb = 6'b101000;
 17'b00000011111000010 : data_comb = 6'b111000;
 17'b00000011111000011 : data_comb = 6'b111000;
 17'b00000011111000100 : data_comb = 6'b111000;
 17'b00000011111000101 : data_comb = 6'b111000;
 17'b00000011111000110 : data_comb = 6'b111000;
 17'b00000011111000111 : data_comb = 6'b111000;
 17'b00000011111001000 : data_comb = 6'b111000;
 17'b00000011111001001 : data_comb = 6'b111000;
 17'b00000011111001010 : data_comb = 6'b111000;
 17'b00000011111001011 : data_comb = 6'b111000;
 17'b00000011111001100 : data_comb = 6'b010101;
 17'b00000011111001101 : data_comb = 6'b000101;
 17'b00000011111001110 : data_comb = 6'b000101;
 17'b00000011111001111 : data_comb = 6'b000101;
 17'b00000011111010000 : data_comb = 6'b000101;
 17'b00000011111010001 : data_comb = 6'b000101;
 17'b00000011111010010 : data_comb = 6'b010101;
 17'b00000011111010011 : data_comb = 6'b111000;
 17'b00000011111010100 : data_comb = 6'b111000;
 17'b00000011111010101 : data_comb = 6'b111000;
 17'b00000011111010110 : data_comb = 6'b101000;
 17'b00000011111010111 : data_comb = 6'b111000;
 17'b00000011111011000 : data_comb = 6'b111000;
 17'b00000011111011001 : data_comb = 6'b111000;
 17'b00000011111011010 : data_comb = 6'b111000;
 17'b00000011111011011 : data_comb = 6'b111000;
 17'b00000011111011100 : data_comb = 6'b010101;
 17'b00000011111011101 : data_comb = 6'b000101;
 17'b00000011111011110 : data_comb = 6'b000101;
 17'b00000011111011111 : data_comb = 6'b000101;
 17'b00000011111100000 : data_comb = 6'b000101;
 17'b00000011111100001 : data_comb = 6'b000101;
 17'b00000011111100010 : data_comb = 6'b000101;
 17'b00000011111100011 : data_comb = 6'b000101;
 17'b00000011111100100 : data_comb = 6'b000101;
 17'b00000011111100101 : data_comb = 6'b000101;
 17'b00000011111100110 : data_comb = 6'b000101;
 17'b00000011111100111 : data_comb = 6'b000101;
 17'b00000011111101000 : data_comb = 6'b000101;
 17'b00000011111101001 : data_comb = 6'b000101;
 17'b00000011111101010 : data_comb = 6'b000101;
 17'b00000011111101011 : data_comb = 6'b000101;
 17'b00000011111101100 : data_comb = 6'b000101;
 17'b00000011111101101 : data_comb = 6'b000101;
 17'b00000011111101110 : data_comb = 6'b000101;
 17'b00000011111101111 : data_comb = 6'b000101;
 17'b00000011111110000 : data_comb = 6'b000101;
 17'b00000011111110001 : data_comb = 6'b000101;
 17'b00000011111110010 : data_comb = 6'b000101;
 17'b00000011111110011 : data_comb = 6'b000101;
 17'b00000011111110100 : data_comb = 6'b000101;
 17'b00000011111110101 : data_comb = 6'b000101;
 17'b00000011111110110 : data_comb = 6'b000101;
 17'b00000011111110111 : data_comb = 6'b000101;
 17'b00000011111111000 : data_comb = 6'b000101;
 17'b00000011111111001 : data_comb = 6'b000101;
 17'b00000011111111010 : data_comb = 6'b000101;
 17'b00000011111111011 : data_comb = 6'b000101;
 17'b00000011111111100 : data_comb = 6'b000101;
 17'b00000011111111101 : data_comb = 6'b000101;
 17'b00000011111111110 : data_comb = 6'b000101;
 17'b00000011111111111 : data_comb = 6'b000101;
 17'b00000100000000000 : data_comb = 6'b000101;
 17'b00000100000000001 : data_comb = 6'b000101;
 17'b00000100000000010 : data_comb = 6'b000101;
 17'b00000100000000011 : data_comb = 6'b000101;
 17'b00000100000000100 : data_comb = 6'b000101;
 17'b00000100000000101 : data_comb = 6'b000101;
 17'b00000100000000110 : data_comb = 6'b000101;
 17'b00000100000000111 : data_comb = 6'b000101;
 17'b00000100000001000 : data_comb = 6'b000101;
 17'b00000100000001001 : data_comb = 6'b000101;
 17'b00000100000001010 : data_comb = 6'b000101;
 17'b00000100000001011 : data_comb = 6'b000101;
 17'b00000100000001100 : data_comb = 6'b000101;
 17'b00000100000001101 : data_comb = 6'b000101;
 17'b00000100000001110 : data_comb = 6'b000101;
 17'b00000100000001111 : data_comb = 6'b000101;
 17'b00000100000010000 : data_comb = 6'b000101;
 17'b00000100000010001 : data_comb = 6'b010101;
 17'b00000100000010010 : data_comb = 6'b111000;
 17'b00000100000010011 : data_comb = 6'b111000;
 17'b00000100000010100 : data_comb = 6'b111000;
 17'b00000100000010101 : data_comb = 6'b111000;
 17'b00000100000010110 : data_comb = 6'b111000;
 17'b00000100000010111 : data_comb = 6'b111000;
 17'b00000100000011000 : data_comb = 6'b111000;
 17'b00000100000011001 : data_comb = 6'b111000;
 17'b00000100000011010 : data_comb = 6'b111000;
 17'b00000100000011011 : data_comb = 6'b111000;
 17'b00000100000011100 : data_comb = 6'b101000;
 17'b00000100000011101 : data_comb = 6'b101000;
 17'b00000100000011110 : data_comb = 6'b000101;
 17'b00000100000011111 : data_comb = 6'b000101;
 17'b00000100000100000 : data_comb = 6'b000101;
 17'b00000100000100001 : data_comb = 6'b000110;
 17'b00000100000100010 : data_comb = 6'b101000;
 17'b00000100000100011 : data_comb = 6'b111000;
 17'b00000100000100100 : data_comb = 6'b111000;
 17'b00000100000100101 : data_comb = 6'b111000;
 17'b00000100000100110 : data_comb = 6'b111000;
 17'b00000100000100111 : data_comb = 6'b111000;
 17'b00000100000101000 : data_comb = 6'b111000;
 17'b00000100000101001 : data_comb = 6'b111000;
 17'b00000100000101010 : data_comb = 6'b111000;
 17'b00000100000101011 : data_comb = 6'b101000;
 17'b00000100000101100 : data_comb = 6'b000101;
 17'b00000100000101101 : data_comb = 6'b000101;
 17'b00000100000101110 : data_comb = 6'b000101;
 17'b00000100000101111 : data_comb = 6'b011001;
 17'b00000100000110000 : data_comb = 6'b011001;
 17'b00000100000110001 : data_comb = 6'b011001;
 17'b00000100000110010 : data_comb = 6'b011001;
 17'b00000100000110011 : data_comb = 6'b011001;
 17'b00000100000110100 : data_comb = 6'b011001;
 17'b00000100000110101 : data_comb = 6'b011001;
 17'b00000100000110110 : data_comb = 6'b011001;
 17'b00000100000110111 : data_comb = 6'b011001;
 17'b00000100000111000 : data_comb = 6'b011001;
 17'b00000100000111001 : data_comb = 6'b011001;
 17'b00000100000111010 : data_comb = 6'b011001;
 17'b00000100000111011 : data_comb = 6'b011001;
 17'b00000100000111100 : data_comb = 6'b000101;
 17'b00000100000111101 : data_comb = 6'b000101;
 17'b00000100000111110 : data_comb = 6'b000101;
 17'b00000100000111111 : data_comb = 6'b000101;
 17'b00000100001000000 : data_comb = 6'b000101;
 17'b00000100001000001 : data_comb = 6'b000101;
 17'b00000100001000010 : data_comb = 6'b000101;
 17'b00000100001000011 : data_comb = 6'b000101;
 17'b00000100001000100 : data_comb = 6'b000101;
 17'b00000100001000101 : data_comb = 6'b000101;
 17'b00000100001000110 : data_comb = 6'b000101;
 17'b00000100001000111 : data_comb = 6'b000101;
 17'b00000100001001000 : data_comb = 6'b000101;
 17'b00000100001001001 : data_comb = 6'b000101;
 17'b00000100001001010 : data_comb = 6'b000101;
 17'b00000100001001011 : data_comb = 6'b010101;
 17'b00000100001001100 : data_comb = 6'b100101;
 17'b00000100001001101 : data_comb = 6'b010101;
 17'b00000100001001110 : data_comb = 6'b000101;
 17'b00000100001001111 : data_comb = 6'b000101;
 17'b00000100001010000 : data_comb = 6'b000101;
 17'b00000100001010001 : data_comb = 6'b000101;
 17'b00000100001010010 : data_comb = 6'b000101;
 17'b00000100001010011 : data_comb = 6'b000101;
 17'b00000100001010100 : data_comb = 6'b011001;
 17'b00000100001010101 : data_comb = 6'b011001;
 17'b00000100001010110 : data_comb = 6'b011001;
 17'b00000100001010111 : data_comb = 6'b011001;
 17'b00000100001011000 : data_comb = 6'b011001;
 17'b00000100001011001 : data_comb = 6'b011001;
 17'b00000100001011010 : data_comb = 6'b011001;
 17'b00000100001011011 : data_comb = 6'b011001;
 17'b00000100001011100 : data_comb = 6'b011001;
 17'b00000100001011101 : data_comb = 6'b011001;
 17'b00000100001011110 : data_comb = 6'b011001;
 17'b00000100001011111 : data_comb = 6'b011001;
 17'b00000100001100000 : data_comb = 6'b001001;
 17'b00000100001100001 : data_comb = 6'b011001;
 17'b00000100001100010 : data_comb = 6'b111000;
 17'b00000100001100011 : data_comb = 6'b111000;
 17'b00000100001100100 : data_comb = 6'b111000;
 17'b00000100001100101 : data_comb = 6'b111000;
 17'b00000100001100110 : data_comb = 6'b111000;
 17'b00000100001100111 : data_comb = 6'b111000;
 17'b00000100001101000 : data_comb = 6'b111000;
 17'b00000100001101001 : data_comb = 6'b111000;
 17'b00000100001101010 : data_comb = 6'b111000;
 17'b00000100001101011 : data_comb = 6'b101000;
 17'b00000100001101100 : data_comb = 6'b101000;
 17'b00000100001101101 : data_comb = 6'b010101;
 17'b00000100001101110 : data_comb = 6'b000101;
 17'b00000100001101111 : data_comb = 6'b000101;
 17'b00000100001110000 : data_comb = 6'b101001;
 17'b00000100001110001 : data_comb = 6'b111000;
 17'b00000100001110010 : data_comb = 6'b111000;
 17'b00000100001110011 : data_comb = 6'b111000;
 17'b00000100001110100 : data_comb = 6'b111000;
 17'b00000100001110101 : data_comb = 6'b111000;
 17'b00000100001110110 : data_comb = 6'b111000;
 17'b00000100001110111 : data_comb = 6'b111000;
 17'b00000100001111000 : data_comb = 6'b111000;
 17'b00000100001111001 : data_comb = 6'b111000;
 17'b00000100001111010 : data_comb = 6'b111000;
 17'b00000100001111011 : data_comb = 6'b011001;
 17'b00000100001111100 : data_comb = 6'b010101;
 17'b00000100001111101 : data_comb = 6'b000101;
 17'b00000100001111110 : data_comb = 6'b000101;
 17'b00000100001111111 : data_comb = 6'b011000;
 17'b00000100010000000 : data_comb = 6'b011000;
 17'b00000100010000001 : data_comb = 6'b011000;
 17'b00000100010000010 : data_comb = 6'b011000;
 17'b00000100010000011 : data_comb = 6'b011000;
 17'b00000100010000100 : data_comb = 6'b011000;
 17'b00000100010000101 : data_comb = 6'b011000;
 17'b00000100010000110 : data_comb = 6'b011000;
 17'b00000100010000111 : data_comb = 6'b011000;
 17'b00000100010001000 : data_comb = 6'b011000;
 17'b00000100010001001 : data_comb = 6'b011000;
 17'b00000100010001010 : data_comb = 6'b011000;
 17'b00000100010001011 : data_comb = 6'b011000;
 17'b00000100010001100 : data_comb = 6'b011000;
 17'b00000100010001101 : data_comb = 6'b000101;
 17'b00000100010001110 : data_comb = 6'b000101;
 17'b00000100010001111 : data_comb = 6'b000101;
 17'b00000100010010000 : data_comb = 6'b000101;
 17'b00000100010010001 : data_comb = 6'b000101;
 17'b00000100010010010 : data_comb = 6'b000101;
 17'b00000100010010011 : data_comb = 6'b000101;
 17'b00000100010010100 : data_comb = 6'b000101;
 17'b00000100010010101 : data_comb = 6'b000101;
 17'b00000100010010110 : data_comb = 6'b000101;
 17'b00000100010010111 : data_comb = 6'b000101;
 17'b00000100010011000 : data_comb = 6'b000101;
 17'b00000100010011001 : data_comb = 6'b000101;
 17'b00000100010011010 : data_comb = 6'b101000;
 17'b00000100010011011 : data_comb = 6'b111000;
 17'b00000100010011100 : data_comb = 6'b111000;
 17'b00000100010011101 : data_comb = 6'b111000;
 17'b00000100010011110 : data_comb = 6'b010101;
 17'b00000100010011111 : data_comb = 6'b000101;
 17'b00000100010100000 : data_comb = 6'b000101;
 17'b00000100010100001 : data_comb = 6'b000101;
 17'b00000100010100010 : data_comb = 6'b000101;
 17'b00000100010100011 : data_comb = 6'b000101;
 17'b00000100010100100 : data_comb = 6'b011000;
 17'b00000100010100101 : data_comb = 6'b011000;
 17'b00000100010100110 : data_comb = 6'b011000;
 17'b00000100010100111 : data_comb = 6'b011000;
 17'b00000100010101000 : data_comb = 6'b011000;
 17'b00000100010101001 : data_comb = 6'b011000;
 17'b00000100010101010 : data_comb = 6'b011000;
 17'b00000100010101011 : data_comb = 6'b011000;
 17'b00000100010101100 : data_comb = 6'b011000;
 17'b00000100010101101 : data_comb = 6'b011000;
 17'b00000100010101110 : data_comb = 6'b011000;
 17'b00000100010101111 : data_comb = 6'b011000;
 17'b00000100010110000 : data_comb = 6'b011000;
 17'b00000100010110001 : data_comb = 6'b011000;
 17'b00000100010110010 : data_comb = 6'b111000;
 17'b00000100010110011 : data_comb = 6'b111000;
 17'b00000100010110100 : data_comb = 6'b111000;
 17'b00000100010110101 : data_comb = 6'b111000;
 17'b00000100010110110 : data_comb = 6'b111000;
 17'b00000100010110111 : data_comb = 6'b111000;
 17'b00000100010111000 : data_comb = 6'b010101;
 17'b00000100010111001 : data_comb = 6'b000101;
 17'b00000100010111010 : data_comb = 6'b000101;
 17'b00000100010111011 : data_comb = 6'b000101;
 17'b00000100010111100 : data_comb = 6'b000101;
 17'b00000100010111101 : data_comb = 6'b000101;
 17'b00000100010111110 : data_comb = 6'b000101;
 17'b00000100010111111 : data_comb = 6'b000101;
 17'b00000100011000000 : data_comb = 6'b111000;
 17'b00000100011000001 : data_comb = 6'b111000;
 17'b00000100011000010 : data_comb = 6'b111000;
 17'b00000100011000011 : data_comb = 6'b111000;
 17'b00000100011000100 : data_comb = 6'b111000;
 17'b00000100011000101 : data_comb = 6'b111000;
 17'b00000100011000110 : data_comb = 6'b111000;
 17'b00000100011000111 : data_comb = 6'b111000;
 17'b00000100011001000 : data_comb = 6'b111000;
 17'b00000100011001001 : data_comb = 6'b111000;
 17'b00000100011001010 : data_comb = 6'b111000;
 17'b00000100011001011 : data_comb = 6'b111000;
 17'b00000100011001100 : data_comb = 6'b111000;
 17'b00000100011001101 : data_comb = 6'b000101;
 17'b00000100011001110 : data_comb = 6'b000101;
 17'b00000100011001111 : data_comb = 6'b000100;
 17'b00000100011010000 : data_comb = 6'b011000;
 17'b00000100011010001 : data_comb = 6'b000100;
 17'b00000100011010010 : data_comb = 6'b010100;
 17'b00000100011010011 : data_comb = 6'b011000;
 17'b00000100011010100 : data_comb = 6'b011000;
 17'b00000100011010101 : data_comb = 6'b000100;
 17'b00000100011010110 : data_comb = 6'b010100;
 17'b00000100011010111 : data_comb = 6'b011000;
 17'b00000100011011000 : data_comb = 6'b011000;
 17'b00000100011011001 : data_comb = 6'b000100;
 17'b00000100011011010 : data_comb = 6'b010100;
 17'b00000100011011011 : data_comb = 6'b011000;
 17'b00000100011011100 : data_comb = 6'b000101;
 17'b00000100011011101 : data_comb = 6'b000101;
 17'b00000100011011110 : data_comb = 6'b000101;
 17'b00000100011011111 : data_comb = 6'b000101;
 17'b00000100011100000 : data_comb = 6'b000101;
 17'b00000100011100001 : data_comb = 6'b000101;
 17'b00000100011100010 : data_comb = 6'b000101;
 17'b00000100011100011 : data_comb = 6'b000101;
 17'b00000100011100100 : data_comb = 6'b000101;
 17'b00000100011100101 : data_comb = 6'b000101;
 17'b00000100011100110 : data_comb = 6'b000101;
 17'b00000100011100111 : data_comb = 6'b000101;
 17'b00000100011101000 : data_comb = 6'b000101;
 17'b00000100011101001 : data_comb = 6'b000101;
 17'b00000100011101010 : data_comb = 6'b111000;
 17'b00000100011101011 : data_comb = 6'b111000;
 17'b00000100011101100 : data_comb = 6'b111000;
 17'b00000100011101101 : data_comb = 6'b111000;
 17'b00000100011101110 : data_comb = 6'b111000;
 17'b00000100011101111 : data_comb = 6'b000101;
 17'b00000100011110000 : data_comb = 6'b000101;
 17'b00000100011110001 : data_comb = 6'b000101;
 17'b00000100011110010 : data_comb = 6'b000101;
 17'b00000100011110011 : data_comb = 6'b000101;
 17'b00000100011110100 : data_comb = 6'b000100;
 17'b00000100011110101 : data_comb = 6'b011000;
 17'b00000100011110110 : data_comb = 6'b000100;
 17'b00000100011110111 : data_comb = 6'b010100;
 17'b00000100011111000 : data_comb = 6'b011000;
 17'b00000100011111001 : data_comb = 6'b011000;
 17'b00000100011111010 : data_comb = 6'b000100;
 17'b00000100011111011 : data_comb = 6'b010100;
 17'b00000100011111100 : data_comb = 6'b011000;
 17'b00000100011111101 : data_comb = 6'b011000;
 17'b00000100011111110 : data_comb = 6'b000100;
 17'b00000100011111111 : data_comb = 6'b010100;
 17'b00000100100000000 : data_comb = 6'b011000;
 17'b00000100100000001 : data_comb = 6'b010100;
 17'b00000100100000010 : data_comb = 6'b111000;
 17'b00000100100000011 : data_comb = 6'b111000;
 17'b00000100100000100 : data_comb = 6'b111000;
 17'b00000100100000101 : data_comb = 6'b111000;
 17'b00000100100000110 : data_comb = 6'b111000;
 17'b00000100100000111 : data_comb = 6'b101000;
 17'b00000100100001000 : data_comb = 6'b000101;
 17'b00000100100001001 : data_comb = 6'b000101;
 17'b00000100100001010 : data_comb = 6'b000101;
 17'b00000100100001011 : data_comb = 6'b000101;
 17'b00000100100001100 : data_comb = 6'b000101;
 17'b00000100100001101 : data_comb = 6'b000101;
 17'b00000100100001110 : data_comb = 6'b000101;
 17'b00000100100001111 : data_comb = 6'b000101;
 17'b00000100100010000 : data_comb = 6'b111000;
 17'b00000100100010001 : data_comb = 6'b111000;
 17'b00000100100010010 : data_comb = 6'b111000;
 17'b00000100100010011 : data_comb = 6'b111000;
 17'b00000100100010100 : data_comb = 6'b111000;
 17'b00000100100010101 : data_comb = 6'b111000;
 17'b00000100100010110 : data_comb = 6'b111000;
 17'b00000100100010111 : data_comb = 6'b111000;
 17'b00000100100011000 : data_comb = 6'b111000;
 17'b00000100100011001 : data_comb = 6'b111000;
 17'b00000100100011010 : data_comb = 6'b111000;
 17'b00000100100011011 : data_comb = 6'b111000;
 17'b00000100100011100 : data_comb = 6'b111000;
 17'b00000100100011101 : data_comb = 6'b111000;
 17'b00000100100011110 : data_comb = 6'b000101;
 17'b00000100100011111 : data_comb = 6'b000100;
 17'b00000100100100000 : data_comb = 6'b000100;
 17'b00000100100100001 : data_comb = 6'b000000;
 17'b00000100100100010 : data_comb = 6'b000000;
 17'b00000100100100011 : data_comb = 6'b010100;
 17'b00000100100100100 : data_comb = 6'b000100;
 17'b00000100100100101 : data_comb = 6'b000000;
 17'b00000100100100110 : data_comb = 6'b000000;
 17'b00000100100100111 : data_comb = 6'b000100;
 17'b00000100100101000 : data_comb = 6'b000100;
 17'b00000100100101001 : data_comb = 6'b000000;
 17'b00000100100101010 : data_comb = 6'b000000;
 17'b00000100100101011 : data_comb = 6'b000100;
 17'b00000100100101100 : data_comb = 6'b000101;
 17'b00000100100101101 : data_comb = 6'b000101;
 17'b00000100100101110 : data_comb = 6'b000101;
 17'b00000100100101111 : data_comb = 6'b000101;
 17'b00000100100110000 : data_comb = 6'b000101;
 17'b00000100100110001 : data_comb = 6'b000101;
 17'b00000100100110010 : data_comb = 6'b000101;
 17'b00000100100110011 : data_comb = 6'b000101;
 17'b00000100100110100 : data_comb = 6'b000101;
 17'b00000100100110101 : data_comb = 6'b000101;
 17'b00000100100110110 : data_comb = 6'b000101;
 17'b00000100100110111 : data_comb = 6'b000101;
 17'b00000100100111000 : data_comb = 6'b101000;
 17'b00000100100111001 : data_comb = 6'b111000;
 17'b00000100100111010 : data_comb = 6'b111000;
 17'b00000100100111011 : data_comb = 6'b111000;
 17'b00000100100111100 : data_comb = 6'b111000;
 17'b00000100100111101 : data_comb = 6'b111000;
 17'b00000100100111110 : data_comb = 6'b111000;
 17'b00000100100111111 : data_comb = 6'b111000;
 17'b00000100101000000 : data_comb = 6'b111000;
 17'b00000100101000001 : data_comb = 6'b000101;
 17'b00000100101000010 : data_comb = 6'b000101;
 17'b00000100101000011 : data_comb = 6'b000101;
 17'b00000100101000100 : data_comb = 6'b000100;
 17'b00000100101000101 : data_comb = 6'b000100;
 17'b00000100101000110 : data_comb = 6'b000000;
 17'b00000100101000111 : data_comb = 6'b000000;
 17'b00000100101001000 : data_comb = 6'b010100;
 17'b00000100101001001 : data_comb = 6'b000100;
 17'b00000100101001010 : data_comb = 6'b000000;
 17'b00000100101001011 : data_comb = 6'b000000;
 17'b00000100101001100 : data_comb = 6'b010100;
 17'b00000100101001101 : data_comb = 6'b010100;
 17'b00000100101001110 : data_comb = 6'b000000;
 17'b00000100101001111 : data_comb = 6'b000000;
 17'b00000100101010000 : data_comb = 6'b000100;
 17'b00000100101010001 : data_comb = 6'b010100;
 17'b00000100101010010 : data_comb = 6'b111000;
 17'b00000100101010011 : data_comb = 6'b111000;
 17'b00000100101010100 : data_comb = 6'b111000;
 17'b00000100101010101 : data_comb = 6'b111000;
 17'b00000100101010110 : data_comb = 6'b111000;
 17'b00000100101010111 : data_comb = 6'b111000;
 17'b00000100101011000 : data_comb = 6'b111000;
 17'b00000100101011001 : data_comb = 6'b111000;
 17'b00000100101011010 : data_comb = 6'b111000;
 17'b00000100101011011 : data_comb = 6'b010101;
 17'b00000100101011100 : data_comb = 6'b000101;
 17'b00000100101011101 : data_comb = 6'b000101;
 17'b00000100101011110 : data_comb = 6'b000101;
 17'b00000100101011111 : data_comb = 6'b000101;
 17'b00000100101100000 : data_comb = 6'b010101;
 17'b00000100101100001 : data_comb = 6'b010101;
 17'b00000100101100010 : data_comb = 6'b010101;
 17'b00000100101100011 : data_comb = 6'b010101;
 17'b00000100101100100 : data_comb = 6'b010101;
 17'b00000100101100101 : data_comb = 6'b101001;
 17'b00000100101100110 : data_comb = 6'b111000;
 17'b00000100101100111 : data_comb = 6'b111000;
 17'b00000100101101000 : data_comb = 6'b111000;
 17'b00000100101101001 : data_comb = 6'b111000;
 17'b00000100101101010 : data_comb = 6'b111000;
 17'b00000100101101011 : data_comb = 6'b111000;
 17'b00000100101101100 : data_comb = 6'b111000;
 17'b00000100101101101 : data_comb = 6'b111000;
 17'b00000100101101110 : data_comb = 6'b000101;
 17'b00000100101101111 : data_comb = 6'b000101;
 17'b00000100101110000 : data_comb = 6'b000000;
 17'b00000100101110001 : data_comb = 6'b000000;
 17'b00000100101110010 : data_comb = 6'b000000;
 17'b00000100101110011 : data_comb = 6'b010000;
 17'b00000100101110100 : data_comb = 6'b000000;
 17'b00000100101110101 : data_comb = 6'b000000;
 17'b00000100101110110 : data_comb = 6'b010000;
 17'b00000100101110111 : data_comb = 6'b010000;
 17'b00000100101111000 : data_comb = 6'b010000;
 17'b00000100101111001 : data_comb = 6'b000000;
 17'b00000100101111010 : data_comb = 6'b000000;
 17'b00000100101111011 : data_comb = 6'b000001;
 17'b00000100101111100 : data_comb = 6'b000101;
 17'b00000100101111101 : data_comb = 6'b000101;
 17'b00000100101111110 : data_comb = 6'b000101;
 17'b00000100101111111 : data_comb = 6'b000101;
 17'b00000100110000000 : data_comb = 6'b000101;
 17'b00000100110000001 : data_comb = 6'b000101;
 17'b00000100110000010 : data_comb = 6'b000101;
 17'b00000100110000011 : data_comb = 6'b000101;
 17'b00000100110000100 : data_comb = 6'b000101;
 17'b00000100110000101 : data_comb = 6'b000101;
 17'b00000100110000110 : data_comb = 6'b000101;
 17'b00000100110000111 : data_comb = 6'b000101;
 17'b00000100110001000 : data_comb = 6'b000101;
 17'b00000100110001001 : data_comb = 6'b000101;
 17'b00000100110001010 : data_comb = 6'b000101;
 17'b00000100110001011 : data_comb = 6'b000101;
 17'b00000100110001100 : data_comb = 6'b000101;
 17'b00000100110001101 : data_comb = 6'b000101;
 17'b00000100110001110 : data_comb = 6'b000101;
 17'b00000100110001111 : data_comb = 6'b000101;
 17'b00000100110010000 : data_comb = 6'b000101;
 17'b00000100110010001 : data_comb = 6'b000101;
 17'b00000100110010010 : data_comb = 6'b000101;
 17'b00000100110010011 : data_comb = 6'b000101;
 17'b00000100110010100 : data_comb = 6'b000101;
 17'b00000100110010101 : data_comb = 6'b000000;
 17'b00000100110010110 : data_comb = 6'b000000;
 17'b00000100110010111 : data_comb = 6'b000000;
 17'b00000100110011000 : data_comb = 6'b010000;
 17'b00000100110011001 : data_comb = 6'b010000;
 17'b00000100110011010 : data_comb = 6'b000000;
 17'b00000100110011011 : data_comb = 6'b000000;
 17'b00000100110011100 : data_comb = 6'b010000;
 17'b00000100110011101 : data_comb = 6'b010000;
 17'b00000100110011110 : data_comb = 6'b000000;
 17'b00000100110011111 : data_comb = 6'b000000;
 17'b00000100110100000 : data_comb = 6'b010000;
 17'b00000100110100001 : data_comb = 6'b111000;
 17'b00000100110100010 : data_comb = 6'b111000;
 17'b00000100110100011 : data_comb = 6'b111000;
 17'b00000100110100100 : data_comb = 6'b111000;
 17'b00000100110100101 : data_comb = 6'b111000;
 17'b00000100110100110 : data_comb = 6'b111000;
 17'b00000100110100111 : data_comb = 6'b111000;
 17'b00000100110101000 : data_comb = 6'b111000;
 17'b00000100110101001 : data_comb = 6'b111000;
 17'b00000100110101010 : data_comb = 6'b111000;
 17'b00000100110101011 : data_comb = 6'b111000;
 17'b00000100110101100 : data_comb = 6'b111000;
 17'b00000100110101101 : data_comb = 6'b010101;
 17'b00000100110101110 : data_comb = 6'b000101;
 17'b00000100110101111 : data_comb = 6'b000101;
 17'b00000100110110000 : data_comb = 6'b000101;
 17'b00000100110110001 : data_comb = 6'b000101;
 17'b00000100110110010 : data_comb = 6'b000101;
 17'b00000100110110011 : data_comb = 6'b000101;
 17'b00000100110110100 : data_comb = 6'b000101;
 17'b00000100110110101 : data_comb = 6'b000101;
 17'b00000100110110110 : data_comb = 6'b101000;
 17'b00000100110110111 : data_comb = 6'b111000;
 17'b00000100110111000 : data_comb = 6'b111000;
 17'b00000100110111001 : data_comb = 6'b111000;
 17'b00000100110111010 : data_comb = 6'b111000;
 17'b00000100110111011 : data_comb = 6'b111000;
 17'b00000100110111100 : data_comb = 6'b111000;
 17'b00000100110111101 : data_comb = 6'b011001;
 17'b00000100110111110 : data_comb = 6'b000101;
 17'b00000100110111111 : data_comb = 6'b000101;
 17'b00000100111000000 : data_comb = 6'b000001;
 17'b00000100111000001 : data_comb = 6'b000000;
 17'b00000100111000010 : data_comb = 6'b010000;
 17'b00000100111000011 : data_comb = 6'b010000;
 17'b00000100111000100 : data_comb = 6'b010000;
 17'b00000100111000101 : data_comb = 6'b000000;
 17'b00000100111000110 : data_comb = 6'b010000;
 17'b00000100111000111 : data_comb = 6'b010000;
 17'b00000100111001000 : data_comb = 6'b010000;
 17'b00000100111001001 : data_comb = 6'b000000;
 17'b00000100111001010 : data_comb = 6'b000000;
 17'b00000100111001011 : data_comb = 6'b000101;
 17'b00000100111001100 : data_comb = 6'b000101;
 17'b00000100111001101 : data_comb = 6'b000101;
 17'b00000100111001110 : data_comb = 6'b000101;
 17'b00000100111001111 : data_comb = 6'b000101;
 17'b00000100111010000 : data_comb = 6'b000101;
 17'b00000100111010001 : data_comb = 6'b000101;
 17'b00000100111010010 : data_comb = 6'b000101;
 17'b00000100111010011 : data_comb = 6'b000101;
 17'b00000100111010100 : data_comb = 6'b000101;
 17'b00000100111010101 : data_comb = 6'b000101;
 17'b00000100111010110 : data_comb = 6'b000101;
 17'b00000100111010111 : data_comb = 6'b000101;
 17'b00000100111011000 : data_comb = 6'b000101;
 17'b00000100111011001 : data_comb = 6'b000101;
 17'b00000100111011010 : data_comb = 6'b000101;
 17'b00000100111011011 : data_comb = 6'b000101;
 17'b00000100111011100 : data_comb = 6'b000101;
 17'b00000100111011101 : data_comb = 6'b000101;
 17'b00000100111011110 : data_comb = 6'b000101;
 17'b00000100111011111 : data_comb = 6'b000101;
 17'b00000100111100000 : data_comb = 6'b000101;
 17'b00000100111100001 : data_comb = 6'b000101;
 17'b00000100111100010 : data_comb = 6'b000101;
 17'b00000100111100011 : data_comb = 6'b000101;
 17'b00000100111100100 : data_comb = 6'b000101;
 17'b00000100111100101 : data_comb = 6'b000101;
 17'b00000100111100110 : data_comb = 6'b000000;
 17'b00000100111100111 : data_comb = 6'b000000;
 17'b00000100111101000 : data_comb = 6'b010000;
 17'b00000100111101001 : data_comb = 6'b010000;
 17'b00000100111101010 : data_comb = 6'b010000;
 17'b00000100111101011 : data_comb = 6'b000000;
 17'b00000100111101100 : data_comb = 6'b010000;
 17'b00000100111101101 : data_comb = 6'b010000;
 17'b00000100111101110 : data_comb = 6'b000000;
 17'b00000100111101111 : data_comb = 6'b000000;
 17'b00000100111110000 : data_comb = 6'b100100;
 17'b00000100111110001 : data_comb = 6'b111000;
 17'b00000100111110010 : data_comb = 6'b111000;
 17'b00000100111110011 : data_comb = 6'b111000;
 17'b00000100111110100 : data_comb = 6'b111000;
 17'b00000100111110101 : data_comb = 6'b111000;
 17'b00000100111110110 : data_comb = 6'b111000;
 17'b00000100111110111 : data_comb = 6'b111000;
 17'b00000100111111000 : data_comb = 6'b111000;
 17'b00000100111111001 : data_comb = 6'b111000;
 17'b00000100111111010 : data_comb = 6'b111000;
 17'b00000100111111011 : data_comb = 6'b111000;
 17'b00000100111111100 : data_comb = 6'b111000;
 17'b00000100111111101 : data_comb = 6'b111000;
 17'b00000100111111110 : data_comb = 6'b010101;
 17'b00000100111111111 : data_comb = 6'b000101;
 17'b00000101000000000 : data_comb = 6'b000101;
 17'b00000101000000001 : data_comb = 6'b000101;
 17'b00000101000000010 : data_comb = 6'b000101;
 17'b00000101000000011 : data_comb = 6'b010101;
 17'b00000101000000100 : data_comb = 6'b010101;
 17'b00000101000000101 : data_comb = 6'b111000;
 17'b00000101000000110 : data_comb = 6'b111000;
 17'b00000101000000111 : data_comb = 6'b111000;
 17'b00000101000001000 : data_comb = 6'b111000;
 17'b00000101000001001 : data_comb = 6'b111000;
 17'b00000101000001010 : data_comb = 6'b111000;
 17'b00000101000001011 : data_comb = 6'b111000;
 17'b00000101000001100 : data_comb = 6'b111000;
 17'b00000101000001101 : data_comb = 6'b111000;
 17'b00000101000001110 : data_comb = 6'b111000;
 17'b00000101000001111 : data_comb = 6'b111000;
 17'b00000101000010000 : data_comb = 6'b111000;
 17'b00000101000010001 : data_comb = 6'b000001;
 17'b00000101000010010 : data_comb = 6'b000001;
 17'b00000101000010011 : data_comb = 6'b000001;
 17'b00000101000010100 : data_comb = 6'b000001;
 17'b00000101000010101 : data_comb = 6'b000001;
 17'b00000101000010110 : data_comb = 6'b000001;
 17'b00000101000010111 : data_comb = 6'b000001;
 17'b00000101000011000 : data_comb = 6'b000001;
 17'b00000101000011001 : data_comb = 6'b000001;
 17'b00000101000011010 : data_comb = 6'b000001;
 17'b00000101000011011 : data_comb = 6'b000101;
 17'b00000101000011100 : data_comb = 6'b000101;
 17'b00000101000011101 : data_comb = 6'b000101;
 17'b00000101000011110 : data_comb = 6'b000101;
 17'b00000101000011111 : data_comb = 6'b000101;
 17'b00000101000100000 : data_comb = 6'b000101;
 17'b00000101000100001 : data_comb = 6'b000101;
 17'b00000101000100010 : data_comb = 6'b000101;
 17'b00000101000100011 : data_comb = 6'b000101;
 17'b00000101000100100 : data_comb = 6'b000101;
 17'b00000101000100101 : data_comb = 6'b000101;
 17'b00000101000100110 : data_comb = 6'b000101;
 17'b00000101000100111 : data_comb = 6'b000101;
 17'b00000101000101000 : data_comb = 6'b000101;
 17'b00000101000101001 : data_comb = 6'b000101;
 17'b00000101000101010 : data_comb = 6'b000101;
 17'b00000101000101011 : data_comb = 6'b000101;
 17'b00000101000101100 : data_comb = 6'b000101;
 17'b00000101000101101 : data_comb = 6'b000101;
 17'b00000101000101110 : data_comb = 6'b000101;
 17'b00000101000101111 : data_comb = 6'b000101;
 17'b00000101000110000 : data_comb = 6'b000101;
 17'b00000101000110001 : data_comb = 6'b000101;
 17'b00000101000110010 : data_comb = 6'b000101;
 17'b00000101000110011 : data_comb = 6'b000101;
 17'b00000101000110100 : data_comb = 6'b000101;
 17'b00000101000110101 : data_comb = 6'b000101;
 17'b00000101000110110 : data_comb = 6'b000001;
 17'b00000101000110111 : data_comb = 6'b000001;
 17'b00000101000111000 : data_comb = 6'b000001;
 17'b00000101000111001 : data_comb = 6'b000001;
 17'b00000101000111010 : data_comb = 6'b000001;
 17'b00000101000111011 : data_comb = 6'b000001;
 17'b00000101000111100 : data_comb = 6'b000001;
 17'b00000101000111101 : data_comb = 6'b010000;
 17'b00000101000111110 : data_comb = 6'b010100;
 17'b00000101000111111 : data_comb = 6'b100100;
 17'b00000101001000000 : data_comb = 6'b111000;
 17'b00000101001000001 : data_comb = 6'b111000;
 17'b00000101001000010 : data_comb = 6'b111000;
 17'b00000101001000011 : data_comb = 6'b111000;
 17'b00000101001000100 : data_comb = 6'b111000;
 17'b00000101001000101 : data_comb = 6'b111000;
 17'b00000101001000110 : data_comb = 6'b111000;
 17'b00000101001000111 : data_comb = 6'b111000;
 17'b00000101001001000 : data_comb = 6'b100101;
 17'b00000101001001001 : data_comb = 6'b000110;
 17'b00000101001001010 : data_comb = 6'b000110;
 17'b00000101001001011 : data_comb = 6'b000101;
 17'b00000101001001100 : data_comb = 6'b000101;
 17'b00000101001001101 : data_comb = 6'b000101;
 17'b00000101001001110 : data_comb = 6'b000101;
 17'b00000101001001111 : data_comb = 6'b000101;
 17'b00000101001010000 : data_comb = 6'b000101;
 17'b00000101001010001 : data_comb = 6'b000101;
 17'b00000101001010010 : data_comb = 6'b101000;
 17'b00000101001010011 : data_comb = 6'b111000;
 17'b00000101001010100 : data_comb = 6'b111000;
 17'b00000101001010101 : data_comb = 6'b111000;
 17'b00000101001010110 : data_comb = 6'b111000;
 17'b00000101001010111 : data_comb = 6'b111000;
 17'b00000101001011000 : data_comb = 6'b111000;
 17'b00000101001011001 : data_comb = 6'b111000;
 17'b00000101001011010 : data_comb = 6'b111000;
 17'b00000101001011011 : data_comb = 6'b111000;
 17'b00000101001011100 : data_comb = 6'b111000;
 17'b00000101001011101 : data_comb = 6'b111000;
 17'b00000101001011110 : data_comb = 6'b111000;
 17'b00000101001011111 : data_comb = 6'b111000;
 17'b00000101001100000 : data_comb = 6'b111000;
 17'b00000101001100001 : data_comb = 6'b101000;
 17'b00000101001100010 : data_comb = 6'b000110;
 17'b00000101001100011 : data_comb = 6'b000101;
 17'b00000101001100100 : data_comb = 6'b000101;
 17'b00000101001100101 : data_comb = 6'b000101;
 17'b00000101001100110 : data_comb = 6'b000101;
 17'b00000101001100111 : data_comb = 6'b000101;
 17'b00000101001101000 : data_comb = 6'b000101;
 17'b00000101001101001 : data_comb = 6'b000101;
 17'b00000101001101010 : data_comb = 6'b000101;
 17'b00000101001101011 : data_comb = 6'b000101;
 17'b00000101001101100 : data_comb = 6'b000101;
 17'b00000101001101101 : data_comb = 6'b000101;
 17'b00000101001101110 : data_comb = 6'b000101;
 17'b00000101001101111 : data_comb = 6'b000101;
 17'b00000101001110000 : data_comb = 6'b000101;
 17'b00000101001110001 : data_comb = 6'b000101;
 17'b00000101001110010 : data_comb = 6'b000101;
 17'b00000101001110011 : data_comb = 6'b000101;
 17'b00000101001110100 : data_comb = 6'b000101;
 17'b00000101001110101 : data_comb = 6'b000101;
 17'b00000101001110110 : data_comb = 6'b000101;
 17'b00000101001110111 : data_comb = 6'b000101;
 17'b00000101001111000 : data_comb = 6'b000101;
 17'b00000101001111001 : data_comb = 6'b000101;
 17'b00000101001111010 : data_comb = 6'b000101;
 17'b00000101001111011 : data_comb = 6'b000101;
 17'b00000101001111100 : data_comb = 6'b000101;
 17'b00000101001111101 : data_comb = 6'b000101;
 17'b00000101001111110 : data_comb = 6'b000101;
 17'b00000101001111111 : data_comb = 6'b000101;
 17'b00000101010000000 : data_comb = 6'b000101;
 17'b00000101010000001 : data_comb = 6'b000101;
 17'b00000101010000010 : data_comb = 6'b000101;
 17'b00000101010000011 : data_comb = 6'b000101;
 17'b00000101010000100 : data_comb = 6'b000101;
 17'b00000101010000101 : data_comb = 6'b000101;
 17'b00000101010000110 : data_comb = 6'b000101;
 17'b00000101010000111 : data_comb = 6'b000101;
 17'b00000101010001000 : data_comb = 6'b000101;
 17'b00000101010001001 : data_comb = 6'b000101;
 17'b00000101010001010 : data_comb = 6'b000110;
 17'b00000101010001011 : data_comb = 6'b000101;
 17'b00000101010001100 : data_comb = 6'b010101;
 17'b00000101010001101 : data_comb = 6'b101000;
 17'b00000101010001110 : data_comb = 6'b111000;
 17'b00000101010001111 : data_comb = 6'b111000;
 17'b00000101010010000 : data_comb = 6'b111000;
 17'b00000101010010001 : data_comb = 6'b111000;
 17'b00000101010010010 : data_comb = 6'b111000;
 17'b00000101010010011 : data_comb = 6'b111000;
 17'b00000101010010100 : data_comb = 6'b101000;
 17'b00000101010010101 : data_comb = 6'b000110;
 17'b00000101010010110 : data_comb = 6'b000110;
 17'b00000101010010111 : data_comb = 6'b000110;
 17'b00000101010011000 : data_comb = 6'b000101;
 17'b00000101010011001 : data_comb = 6'b000101;
 17'b00000101010011010 : data_comb = 6'b000101;
 17'b00000101010011011 : data_comb = 6'b000101;
 17'b00000101010011100 : data_comb = 6'b000101;
 17'b00000101010011101 : data_comb = 6'b000101;
 17'b00000101010011110 : data_comb = 6'b000101;
 17'b00000101010011111 : data_comb = 6'b000101;
 17'b00000101010100000 : data_comb = 6'b000101;
 17'b00000101010100001 : data_comb = 6'b000101;
 17'b00000101010100010 : data_comb = 6'b000101;
 17'b00000101010100011 : data_comb = 6'b000101;
 17'b00000101010100100 : data_comb = 6'b000101;
 17'b00000101010100101 : data_comb = 6'b000101;
 17'b00000101010100110 : data_comb = 6'b000101;
 17'b00000101010100111 : data_comb = 6'b000101;
 17'b00000101010101000 : data_comb = 6'b000101;
 17'b00000101010101001 : data_comb = 6'b010101;
 17'b00000101010101010 : data_comb = 6'b010101;
 17'b00000101010101011 : data_comb = 6'b111000;
 17'b00000101010101100 : data_comb = 6'b111000;
 17'b00000101010101101 : data_comb = 6'b111000;
 17'b00000101010101110 : data_comb = 6'b111000;
 17'b00000101010101111 : data_comb = 6'b111000;
 17'b00000101010110000 : data_comb = 6'b111000;
 17'b00000101010110001 : data_comb = 6'b111000;
 17'b00000101010110010 : data_comb = 6'b101000;
 17'b00000101010110011 : data_comb = 6'b101000;
 17'b00000101010110100 : data_comb = 6'b101000;
 17'b00000101010110101 : data_comb = 6'b000101;
 17'b00000101010110110 : data_comb = 6'b000101;
 17'b00000101010110111 : data_comb = 6'b000101;
 17'b00000101010111000 : data_comb = 6'b000101;
 17'b00000101010111001 : data_comb = 6'b000101;
 17'b00000101010111010 : data_comb = 6'b000101;
 17'b00000101010111011 : data_comb = 6'b000101;
 17'b00000101010111100 : data_comb = 6'b000101;
 17'b00000101010111101 : data_comb = 6'b000101;
 17'b00000101010111110 : data_comb = 6'b000101;
 17'b00000101010111111 : data_comb = 6'b000101;
 17'b00000101011000000 : data_comb = 6'b000101;
 17'b00000101011000001 : data_comb = 6'b000101;
 17'b00000101011000010 : data_comb = 6'b000101;
 17'b00000101011000011 : data_comb = 6'b000101;
 17'b00000101011000100 : data_comb = 6'b000101;
 17'b00000101011000101 : data_comb = 6'b000101;
 17'b00000101011000110 : data_comb = 6'b000101;
 17'b00000101011000111 : data_comb = 6'b000101;
 17'b00000101011001000 : data_comb = 6'b000101;
 17'b00000101011001001 : data_comb = 6'b000101;
 17'b00000101011001010 : data_comb = 6'b000101;
 17'b00000101011001011 : data_comb = 6'b000101;
 17'b00000101011001100 : data_comb = 6'b000101;
 17'b00000101011001101 : data_comb = 6'b000101;
 17'b00000101011001110 : data_comb = 6'b000101;
 17'b00000101011001111 : data_comb = 6'b000101;
 17'b00000101011010000 : data_comb = 6'b000101;
 17'b00000101011010001 : data_comb = 6'b000101;
 17'b00000101011010010 : data_comb = 6'b000101;
 17'b00000101011010011 : data_comb = 6'b000101;
 17'b00000101011010100 : data_comb = 6'b000101;
 17'b00000101011010101 : data_comb = 6'b000101;
 17'b00000101011010110 : data_comb = 6'b000101;
 17'b00000101011010111 : data_comb = 6'b000101;
 17'b00000101011011000 : data_comb = 6'b000101;
 17'b00000101011011001 : data_comb = 6'b010101;
 17'b00000101011011010 : data_comb = 6'b111000;
 17'b00000101011011011 : data_comb = 6'b111000;
 17'b00000101011011100 : data_comb = 6'b111000;
 17'b00000101011011101 : data_comb = 6'b111000;
 17'b00000101011011110 : data_comb = 6'b111000;
 17'b00000101011011111 : data_comb = 6'b111000;
 17'b00000101011100000 : data_comb = 6'b111000;
 17'b00000101011100001 : data_comb = 6'b111000;
 17'b00000101011100010 : data_comb = 6'b111000;
 17'b00000101011100011 : data_comb = 6'b111000;
 17'b00000101011100100 : data_comb = 6'b111000;
 17'b00000101011100101 : data_comb = 6'b101000;
 17'b00000101011100110 : data_comb = 6'b000101;
 17'b00000101011100111 : data_comb = 6'b000101;
 17'b00000101011101000 : data_comb = 6'b000101;
 17'b00000101011101001 : data_comb = 6'b000101;
 17'b00000101011101010 : data_comb = 6'b000101;
 17'b00000101011101011 : data_comb = 6'b000101;
 17'b00000101011101100 : data_comb = 6'b000101;
 17'b00000101011101101 : data_comb = 6'b000101;
 17'b00000101011101110 : data_comb = 6'b000101;
 17'b00000101011101111 : data_comb = 6'b000101;
 17'b00000101011110000 : data_comb = 6'b000110;
 17'b00000101011110001 : data_comb = 6'b000110;
 17'b00000101011110010 : data_comb = 6'b000110;
 17'b00000101011110011 : data_comb = 6'b000110;
 17'b00000101011110100 : data_comb = 6'b000110;
 17'b00000101011110101 : data_comb = 6'b000110;
 17'b00000101011110110 : data_comb = 6'b000110;
 17'b00000101011110111 : data_comb = 6'b000110;
 17'b00000101011111000 : data_comb = 6'b000110;
 17'b00000101011111001 : data_comb = 6'b011001;
 17'b00000101011111010 : data_comb = 6'b111000;
 17'b00000101011111011 : data_comb = 6'b111000;
 17'b00000101011111100 : data_comb = 6'b111000;
 17'b00000101011111101 : data_comb = 6'b111000;
 17'b00000101011111110 : data_comb = 6'b101000;
 17'b00000101011111111 : data_comb = 6'b101001;
 17'b00000101100000000 : data_comb = 6'b101001;
 17'b00000101100000001 : data_comb = 6'b101001;
 17'b00000101100000010 : data_comb = 6'b101001;
 17'b00000101100000011 : data_comb = 6'b101001;
 17'b00000101100000100 : data_comb = 6'b101001;
 17'b00000101100000101 : data_comb = 6'b000110;
 17'b00000101100000110 : data_comb = 6'b000110;
 17'b00000101100000111 : data_comb = 6'b000110;
 17'b00000101100001000 : data_comb = 6'b000110;
 17'b00000101100001001 : data_comb = 6'b000110;
 17'b00000101100001010 : data_comb = 6'b000110;
 17'b00000101100001011 : data_comb = 6'b000110;
 17'b00000101100001100 : data_comb = 6'b000110;
 17'b00000101100001101 : data_comb = 6'b000110;
 17'b00000101100001110 : data_comb = 6'b000110;
 17'b00000101100001111 : data_comb = 6'b000110;
 17'b00000101100010000 : data_comb = 6'b000110;
 17'b00000101100010001 : data_comb = 6'b000110;
 17'b00000101100010010 : data_comb = 6'b000110;
 17'b00000101100010011 : data_comb = 6'b000110;
 17'b00000101100010100 : data_comb = 6'b000110;
 17'b00000101100010101 : data_comb = 6'b000110;
 17'b00000101100010110 : data_comb = 6'b000110;
 17'b00000101100010111 : data_comb = 6'b000110;
 17'b00000101100011000 : data_comb = 6'b000110;
 17'b00000101100011001 : data_comb = 6'b000110;
 17'b00000101100011010 : data_comb = 6'b000110;
 17'b00000101100011011 : data_comb = 6'b000110;
 17'b00000101100011100 : data_comb = 6'b000110;
 17'b00000101100011101 : data_comb = 6'b000110;
 17'b00000101100011110 : data_comb = 6'b000110;
 17'b00000101100011111 : data_comb = 6'b000110;
 17'b00000101100100000 : data_comb = 6'b000110;
 17'b00000101100100001 : data_comb = 6'b000110;
 17'b00000101100100010 : data_comb = 6'b000110;
 17'b00000101100100011 : data_comb = 6'b000110;
 17'b00000101100100100 : data_comb = 6'b101001;
 17'b00000101100100101 : data_comb = 6'b101000;
 17'b00000101100100110 : data_comb = 6'b111000;
 17'b00000101100100111 : data_comb = 6'b111000;
 17'b00000101100101000 : data_comb = 6'b111000;
 17'b00000101100101001 : data_comb = 6'b111000;
 17'b00000101100101010 : data_comb = 6'b111000;
 17'b00000101100101011 : data_comb = 6'b111000;
 17'b00000101100101100 : data_comb = 6'b111000;
 17'b00000101100101101 : data_comb = 6'b111000;
 17'b00000101100101110 : data_comb = 6'b010101;
 17'b00000101100101111 : data_comb = 6'b010101;
 17'b00000101100110000 : data_comb = 6'b010101;
 17'b00000101100110001 : data_comb = 6'b010101;
 17'b00000101100110010 : data_comb = 6'b111000;
 17'b00000101100110011 : data_comb = 6'b111000;
 17'b00000101100110100 : data_comb = 6'b111000;
 17'b00000101100110101 : data_comb = 6'b111000;
 17'b00000101100110110 : data_comb = 6'b010101;
 17'b00000101100110111 : data_comb = 6'b000101;
 17'b00000101100111000 : data_comb = 6'b000101;
 17'b00000101100111001 : data_comb = 6'b000101;
 17'b00000101100111010 : data_comb = 6'b000101;
 17'b00000101100111011 : data_comb = 6'b000101;
 17'b00000101100111100 : data_comb = 6'b000101;
 17'b00000101100111101 : data_comb = 6'b000101;
 17'b00000101100111110 : data_comb = 6'b000101;
 17'b00000101100111111 : data_comb = 6'b000101;
 17'b00000101101000000 : data_comb = 6'b000110;
 17'b00000101101000001 : data_comb = 6'b000110;
 17'b00000101101000010 : data_comb = 6'b000110;
 17'b00000101101000011 : data_comb = 6'b000110;
 17'b00000101101000100 : data_comb = 6'b000110;
 17'b00000101101000101 : data_comb = 6'b000110;
 17'b00000101101000110 : data_comb = 6'b000110;
 17'b00000101101000111 : data_comb = 6'b000110;
 17'b00000101101001000 : data_comb = 6'b000110;
 17'b00000101101001001 : data_comb = 6'b000101;
 17'b00000101101001010 : data_comb = 6'b010101;
 17'b00000101101001011 : data_comb = 6'b010101;
 17'b00000101101001100 : data_comb = 6'b010101;
 17'b00000101101001101 : data_comb = 6'b010101;
 17'b00000101101001110 : data_comb = 6'b000101;
 17'b00000101101001111 : data_comb = 6'b000110;
 17'b00000101101010000 : data_comb = 6'b000110;
 17'b00000101101010001 : data_comb = 6'b000110;
 17'b00000101101010010 : data_comb = 6'b000110;
 17'b00000101101010011 : data_comb = 6'b000110;
 17'b00000101101010100 : data_comb = 6'b000110;
 17'b00000101101010101 : data_comb = 6'b000110;
 17'b00000101101010110 : data_comb = 6'b000110;
 17'b00000101101010111 : data_comb = 6'b000110;
 17'b00000101101011000 : data_comb = 6'b000110;
 17'b00000101101011001 : data_comb = 6'b000110;
 17'b00000101101011010 : data_comb = 6'b000110;
 17'b00000101101011011 : data_comb = 6'b000110;
 17'b00000101101011100 : data_comb = 6'b000110;
 17'b00000101101011101 : data_comb = 6'b000110;
 17'b00000101101011110 : data_comb = 6'b000110;
 17'b00000101101011111 : data_comb = 6'b000110;
 17'b00000101101100000 : data_comb = 6'b000110;
 17'b00000101101100001 : data_comb = 6'b000110;
 17'b00000101101100010 : data_comb = 6'b000110;
 17'b00000101101100011 : data_comb = 6'b000110;
 17'b00000101101100100 : data_comb = 6'b000110;
 17'b00000101101100101 : data_comb = 6'b000110;
 17'b00000101101100110 : data_comb = 6'b000110;
 17'b00000101101100111 : data_comb = 6'b000110;
 17'b00000101101101000 : data_comb = 6'b000110;
 17'b00000101101101001 : data_comb = 6'b000110;
 17'b00000101101101010 : data_comb = 6'b000110;
 17'b00000101101101011 : data_comb = 6'b000110;
 17'b00000101101101100 : data_comb = 6'b000110;
 17'b00000101101101101 : data_comb = 6'b000110;
 17'b00000101101101110 : data_comb = 6'b000110;
 17'b00000101101101111 : data_comb = 6'b000110;
 17'b00000101101110000 : data_comb = 6'b000110;
 17'b00000101101110001 : data_comb = 6'b000110;
 17'b00000101101110010 : data_comb = 6'b000110;
 17'b00000101101110011 : data_comb = 6'b000110;
 17'b00000101101110100 : data_comb = 6'b101000;
 17'b00000101101110101 : data_comb = 6'b101000;
 17'b00000101101110110 : data_comb = 6'b101000;
 17'b00000101101110111 : data_comb = 6'b101000;
 17'b00000101101111000 : data_comb = 6'b101000;
 17'b00000101101111001 : data_comb = 6'b101000;
 17'b00000101101111010 : data_comb = 6'b101000;
 17'b00000101101111011 : data_comb = 6'b101000;
 17'b00000101101111100 : data_comb = 6'b101000;
 17'b00000101101111101 : data_comb = 6'b101001;
 17'b00000101101111110 : data_comb = 6'b000110;
 17'b00000101101111111 : data_comb = 6'b000110;
 17'b00000101110000000 : data_comb = 6'b000110;
 17'b00000101110000001 : data_comb = 6'b000110;
 17'b00000101110000010 : data_comb = 6'b010101;
 17'b00000101110000011 : data_comb = 6'b010101;
 17'b00000101110000100 : data_comb = 6'b010101;
 17'b00000101110000101 : data_comb = 6'b000101;
 17'b00000101110000110 : data_comb = 6'b000101;
 17'b00000101110000111 : data_comb = 6'b000110;
 17'b00000101110001000 : data_comb = 6'b000101;
 17'b00000101110001001 : data_comb = 6'b111000;
 17'b00000101110001010 : data_comb = 6'b111000;
 17'b00000101110001011 : data_comb = 6'b111000;
 17'b00000101110001100 : data_comb = 6'b011001;
 17'b00000101110001101 : data_comb = 6'b000110;
 17'b00000101110001110 : data_comb = 6'b000110;
 17'b00000101110001111 : data_comb = 6'b000110;
 17'b00000101110010000 : data_comb = 6'b000110;
 17'b00000101110010001 : data_comb = 6'b000110;
 17'b00000101110010010 : data_comb = 6'b000110;
 17'b00000101110010011 : data_comb = 6'b000110;
 17'b00000101110010100 : data_comb = 6'b000110;
 17'b00000101110010101 : data_comb = 6'b000110;
 17'b00000101110010110 : data_comb = 6'b000110;
 17'b00000101110010111 : data_comb = 6'b000110;
 17'b00000101110011000 : data_comb = 6'b000110;
 17'b00000101110011001 : data_comb = 6'b000110;
 17'b00000101110011010 : data_comb = 6'b000110;
 17'b00000101110011011 : data_comb = 6'b000110;
 17'b00000101110011100 : data_comb = 6'b000110;
 17'b00000101110011101 : data_comb = 6'b000110;
 17'b00000101110011110 : data_comb = 6'b000110;
 17'b00000101110011111 : data_comb = 6'b000110;
 17'b00000101110100000 : data_comb = 6'b000110;
 17'b00000101110100001 : data_comb = 6'b000110;
 17'b00000101110100010 : data_comb = 6'b000110;
 17'b00000101110100011 : data_comb = 6'b000110;
 17'b00000101110100100 : data_comb = 6'b000110;
 17'b00000101110100101 : data_comb = 6'b000110;
 17'b00000101110100110 : data_comb = 6'b000110;
 17'b00000101110100111 : data_comb = 6'b000110;
 17'b00000101110101000 : data_comb = 6'b000110;
 17'b00000101110101001 : data_comb = 6'b000110;
 17'b00000101110101010 : data_comb = 6'b000110;
 17'b00000101110101011 : data_comb = 6'b000110;
 17'b00000101110101100 : data_comb = 6'b000110;
 17'b00000101110101101 : data_comb = 6'b000110;
 17'b00000101110101110 : data_comb = 6'b000110;
 17'b00000101110101111 : data_comb = 6'b000110;
 17'b00000101110110000 : data_comb = 6'b000110;
 17'b00000101110110001 : data_comb = 6'b000110;
 17'b00000101110110010 : data_comb = 6'b000110;
 17'b00000101110110011 : data_comb = 6'b000110;
 17'b00000101110110100 : data_comb = 6'b000110;
 17'b00000101110110101 : data_comb = 6'b000110;
 17'b00000101110110110 : data_comb = 6'b000110;
 17'b00000101110110111 : data_comb = 6'b000110;
 17'b00000101110111000 : data_comb = 6'b000110;
 17'b00000101110111001 : data_comb = 6'b000110;
 17'b00000101110111010 : data_comb = 6'b000110;
 17'b00000101110111011 : data_comb = 6'b000110;
 17'b00000101110111100 : data_comb = 6'b000110;
 17'b00000101110111101 : data_comb = 6'b000110;
 17'b00000101110111110 : data_comb = 6'b000110;
 17'b00000101110111111 : data_comb = 6'b000110;
 17'b00000101111000000 : data_comb = 6'b000110;
 17'b00000101111000001 : data_comb = 6'b000110;
 17'b00000101111000010 : data_comb = 6'b000110;
 17'b00000101111000011 : data_comb = 6'b000110;
 17'b00000101111000100 : data_comb = 6'b000110;
 17'b00000101111000101 : data_comb = 6'b000110;
 17'b00000101111000110 : data_comb = 6'b000110;
 17'b00000101111000111 : data_comb = 6'b000110;
 17'b00000101111001000 : data_comb = 6'b000110;
 17'b00000101111001001 : data_comb = 6'b000110;
 17'b00000101111001010 : data_comb = 6'b000110;
 17'b00000101111001011 : data_comb = 6'b000110;
 17'b00000101111001100 : data_comb = 6'b000110;
 17'b00000101111001101 : data_comb = 6'b000110;
 17'b00000101111001110 : data_comb = 6'b000110;
 17'b00000101111001111 : data_comb = 6'b000110;
 17'b00000101111010000 : data_comb = 6'b000110;
 17'b00000101111010001 : data_comb = 6'b000110;
 17'b00000101111010010 : data_comb = 6'b000110;
 17'b00000101111010011 : data_comb = 6'b000110;
 17'b00000101111010100 : data_comb = 6'b000110;
 17'b00000101111010101 : data_comb = 6'b000110;
 17'b00000101111010110 : data_comb = 6'b000110;
 17'b00000101111010111 : data_comb = 6'b000110;
 17'b00000101111011000 : data_comb = 6'b101000;
 17'b00000101111011001 : data_comb = 6'b111000;
 17'b00000101111011010 : data_comb = 6'b111000;
 17'b00000101111011011 : data_comb = 6'b111000;
 17'b00000101111011100 : data_comb = 6'b111000;
 17'b00000101111011101 : data_comb = 6'b010101;
 17'b00000101111011110 : data_comb = 6'b000110;
 17'b00000101111011111 : data_comb = 6'b000110;
 17'b00000101111100000 : data_comb = 6'b101000;
 17'b00000101111100001 : data_comb = 6'b000101;
 17'b00000101111100010 : data_comb = 6'b000110;
 17'b00000101111100011 : data_comb = 6'b000110;
 17'b00000101111100100 : data_comb = 6'b000110;
 17'b00000101111100101 : data_comb = 6'b101001;
 17'b00000101111100110 : data_comb = 6'b101000;
 17'b00000101111100111 : data_comb = 6'b011001;
 17'b00000101111101000 : data_comb = 6'b000110;
 17'b00000101111101001 : data_comb = 6'b000110;
 17'b00000101111101010 : data_comb = 6'b000110;
 17'b00000101111101011 : data_comb = 6'b000110;
 17'b00000101111101100 : data_comb = 6'b000110;
 17'b00000101111101101 : data_comb = 6'b000110;
 17'b00000101111101110 : data_comb = 6'b000110;
 17'b00000101111101111 : data_comb = 6'b000110;
 17'b00000101111110000 : data_comb = 6'b000110;
 17'b00000101111110001 : data_comb = 6'b000110;
 17'b00000101111110010 : data_comb = 6'b000110;
 17'b00000101111110011 : data_comb = 6'b000110;
 17'b00000101111110100 : data_comb = 6'b000110;
 17'b00000101111110101 : data_comb = 6'b000110;
 17'b00000101111110110 : data_comb = 6'b000110;
 17'b00000101111110111 : data_comb = 6'b000110;
 17'b00000101111111000 : data_comb = 6'b000110;
 17'b00000101111111001 : data_comb = 6'b000110;
 17'b00000101111111010 : data_comb = 6'b000110;
 17'b00000101111111011 : data_comb = 6'b000110;
 17'b00000101111111100 : data_comb = 6'b000110;
 17'b00000101111111101 : data_comb = 6'b000110;
 17'b00000101111111110 : data_comb = 6'b000110;
 17'b00000101111111111 : data_comb = 6'b000110;
 17'b00000110000000000 : data_comb = 6'b000110;
 17'b00000110000000001 : data_comb = 6'b000110;
 17'b00000110000000010 : data_comb = 6'b000110;
 17'b00000110000000011 : data_comb = 6'b000110;
 17'b00000110000000100 : data_comb = 6'b000110;
 17'b00000110000000101 : data_comb = 6'b000110;
 17'b00000110000000110 : data_comb = 6'b000110;
 17'b00000110000000111 : data_comb = 6'b000110;
 17'b00000110000001000 : data_comb = 6'b000110;
 17'b00000110000001001 : data_comb = 6'b000110;
 17'b00000110000001010 : data_comb = 6'b000110;
 17'b00000110000001011 : data_comb = 6'b000110;
 17'b00000110000001100 : data_comb = 6'b000110;
 17'b00000110000001101 : data_comb = 6'b000110;
 17'b00000110000001110 : data_comb = 6'b000110;
 17'b00000110000001111 : data_comb = 6'b000110;
 17'b00000110000010000 : data_comb = 6'b000110;
 17'b00000110000010001 : data_comb = 6'b000110;
 17'b00000110000010010 : data_comb = 6'b000110;
 17'b00000110000010011 : data_comb = 6'b000110;
 17'b00000110000010100 : data_comb = 6'b000110;
 17'b00000110000010101 : data_comb = 6'b000110;
 17'b00000110000010110 : data_comb = 6'b000110;
 17'b00000110000010111 : data_comb = 6'b000110;
 17'b00000110000011000 : data_comb = 6'b000110;
 17'b00000110000011001 : data_comb = 6'b000110;
 17'b00000110000011010 : data_comb = 6'b000110;
 17'b00000110000011011 : data_comb = 6'b000110;
 17'b00000110000011100 : data_comb = 6'b000110;
 17'b00000110000011101 : data_comb = 6'b000110;
 17'b00000110000011110 : data_comb = 6'b000110;
 17'b00000110000011111 : data_comb = 6'b000110;
 17'b00000110000100000 : data_comb = 6'b000110;
 17'b00000110000100001 : data_comb = 6'b000110;
 17'b00000110000100010 : data_comb = 6'b000110;
 17'b00000110000100011 : data_comb = 6'b000110;
 17'b00000110000100100 : data_comb = 6'b000110;
 17'b00000110000100101 : data_comb = 6'b000110;
 17'b00000110000100110 : data_comb = 6'b000110;
 17'b00000110000100111 : data_comb = 6'b011001;
 17'b00000110000101000 : data_comb = 6'b111000;
 17'b00000110000101001 : data_comb = 6'b111000;
 17'b00000110000101010 : data_comb = 6'b111000;
 17'b00000110000101011 : data_comb = 6'b111000;
 17'b00000110000101100 : data_comb = 6'b111000;
 17'b00000110000101101 : data_comb = 6'b111000;
 17'b00000110000101110 : data_comb = 6'b000101;
 17'b00000110000101111 : data_comb = 6'b000110;
 17'b00000110000110000 : data_comb = 6'b111000;
 17'b00000110000110001 : data_comb = 6'b101000;
 17'b00000110000110010 : data_comb = 6'b000101;
 17'b00000110000110011 : data_comb = 6'b000101;
 17'b00000110000110100 : data_comb = 6'b101000;
 17'b00000110000110101 : data_comb = 6'b111000;
 17'b00000110000110110 : data_comb = 6'b111000;
 17'b00000110000110111 : data_comb = 6'b111000;
 17'b00000110000111000 : data_comb = 6'b111000;
 17'b00000110000111001 : data_comb = 6'b000110;
 17'b00000110000111010 : data_comb = 6'b000110;
 17'b00000110000111011 : data_comb = 6'b000110;
 17'b00000110000111100 : data_comb = 6'b000110;
 17'b00000110000111101 : data_comb = 6'b000110;
 17'b00000110000111110 : data_comb = 6'b000110;
 17'b00000110000111111 : data_comb = 6'b000110;
 17'b00000110001000000 : data_comb = 6'b000110;
 17'b00000110001000001 : data_comb = 6'b000110;
 17'b00000110001000010 : data_comb = 6'b000110;
 17'b00000110001000011 : data_comb = 6'b000110;
 17'b00000110001000100 : data_comb = 6'b000110;
 17'b00000110001000101 : data_comb = 6'b000110;
 17'b00000110001000110 : data_comb = 6'b000110;
 17'b00000110001000111 : data_comb = 6'b000110;
 17'b00000110001001000 : data_comb = 6'b000110;
 17'b00000110001001001 : data_comb = 6'b000110;
 17'b00000110001001010 : data_comb = 6'b000110;
 17'b00000110001001011 : data_comb = 6'b000110;
 17'b00000110001001100 : data_comb = 6'b000110;
 17'b00000110001001101 : data_comb = 6'b000110;
 17'b00000110001001110 : data_comb = 6'b000110;
 17'b00000110001001111 : data_comb = 6'b000110;
 17'b00000110001010000 : data_comb = 6'b000110;
 17'b00000110001010001 : data_comb = 6'b000110;
 17'b00000110001010010 : data_comb = 6'b000110;
 17'b00000110001010011 : data_comb = 6'b000110;
 17'b00000110001010100 : data_comb = 6'b000110;
 17'b00000110001010101 : data_comb = 6'b000110;
 17'b00000110001010110 : data_comb = 6'b000110;
 17'b00000110001010111 : data_comb = 6'b000110;
 17'b00000110001011000 : data_comb = 6'b000110;
 17'b00000110001011001 : data_comb = 6'b000110;
 17'b00000110001011010 : data_comb = 6'b000110;
 17'b00000110001011011 : data_comb = 6'b000110;
 17'b00000110001011100 : data_comb = 6'b000110;
 17'b00000110001011101 : data_comb = 6'b000110;
 17'b00000110001011110 : data_comb = 6'b000110;
 17'b00000110001011111 : data_comb = 6'b000110;
 17'b00000110001100000 : data_comb = 6'b000110;
 17'b00000110001100001 : data_comb = 6'b000110;
 17'b00000110001100010 : data_comb = 6'b000110;
 17'b00000110001100011 : data_comb = 6'b000110;
 17'b00000110001100100 : data_comb = 6'b000110;
 17'b00000110001100101 : data_comb = 6'b000110;
 17'b00000110001100110 : data_comb = 6'b000110;
 17'b00000110001100111 : data_comb = 6'b000110;
 17'b00000110001101000 : data_comb = 6'b000110;
 17'b00000110001101001 : data_comb = 6'b000110;
 17'b00000110001101010 : data_comb = 6'b000110;
 17'b00000110001101011 : data_comb = 6'b000110;
 17'b00000110001101100 : data_comb = 6'b000110;
 17'b00000110001101101 : data_comb = 6'b000110;
 17'b00000110001101110 : data_comb = 6'b000110;
 17'b00000110001101111 : data_comb = 6'b000110;
 17'b00000110001110000 : data_comb = 6'b000110;
 17'b00000110001110001 : data_comb = 6'b000110;
 17'b00000110001110010 : data_comb = 6'b000110;
 17'b00000110001110011 : data_comb = 6'b000110;
 17'b00000110001110100 : data_comb = 6'b000110;
 17'b00000110001110101 : data_comb = 6'b000110;
 17'b00000110001110110 : data_comb = 6'b000110;
 17'b00000110001110111 : data_comb = 6'b111000;
 17'b00000110001111000 : data_comb = 6'b111000;
 17'b00000110001111001 : data_comb = 6'b111000;
 17'b00000110001111010 : data_comb = 6'b111000;
 17'b00000110001111011 : data_comb = 6'b111000;
 17'b00000110001111100 : data_comb = 6'b111000;
 17'b00000110001111101 : data_comb = 6'b111000;
 17'b00000110001111110 : data_comb = 6'b000101;
 17'b00000110001111111 : data_comb = 6'b000110;
 17'b00000110010000000 : data_comb = 6'b111000;
 17'b00000110010000001 : data_comb = 6'b111000;
 17'b00000110010000010 : data_comb = 6'b111000;
 17'b00000110010000011 : data_comb = 6'b101000;
 17'b00000110010000100 : data_comb = 6'b111000;
 17'b00000110010000101 : data_comb = 6'b111000;
 17'b00000110010000110 : data_comb = 6'b111000;
 17'b00000110010000111 : data_comb = 6'b111000;
 17'b00000110010001000 : data_comb = 6'b111000;
 17'b00000110010001001 : data_comb = 6'b000110;
 17'b00000110010001010 : data_comb = 6'b000110;
 17'b00000110010001011 : data_comb = 6'b000110;
 17'b00000110010001100 : data_comb = 6'b000110;
 17'b00000110010001101 : data_comb = 6'b000110;
 17'b00000110010001110 : data_comb = 6'b000110;
 17'b00000110010001111 : data_comb = 6'b000110;
 17'b00000110010010000 : data_comb = 6'b000110;
 17'b00000110010010001 : data_comb = 6'b000101;
 17'b00000110010010010 : data_comb = 6'b000101;
 17'b00000110010010011 : data_comb = 6'b000110;
 17'b00000110010010100 : data_comb = 6'b000110;
 17'b00000110010010101 : data_comb = 6'b000110;
 17'b00000110010010110 : data_comb = 6'b000110;
 17'b00000110010010111 : data_comb = 6'b000110;
 17'b00000110010011000 : data_comb = 6'b000110;
 17'b00000110010011001 : data_comb = 6'b000101;
 17'b00000110010011010 : data_comb = 6'b000101;
 17'b00000110010011011 : data_comb = 6'b000110;
 17'b00000110010011100 : data_comb = 6'b000110;
 17'b00000110010011101 : data_comb = 6'b000110;
 17'b00000110010011110 : data_comb = 6'b000110;
 17'b00000110010011111 : data_comb = 6'b000110;
 17'b00000110010100000 : data_comb = 6'b000110;
 17'b00000110010100001 : data_comb = 6'b000110;
 17'b00000110010100010 : data_comb = 6'b000110;
 17'b00000110010100011 : data_comb = 6'b000110;
 17'b00000110010100100 : data_comb = 6'b000110;
 17'b00000110010100101 : data_comb = 6'b000101;
 17'b00000110010100110 : data_comb = 6'b000101;
 17'b00000110010100111 : data_comb = 6'b000101;
 17'b00000110010101000 : data_comb = 6'b000110;
 17'b00000110010101001 : data_comb = 6'b000110;
 17'b00000110010101010 : data_comb = 6'b000110;
 17'b00000110010101011 : data_comb = 6'b000110;
 17'b00000110010101100 : data_comb = 6'b000110;
 17'b00000110010101101 : data_comb = 6'b000110;
 17'b00000110010101110 : data_comb = 6'b000110;
 17'b00000110010101111 : data_comb = 6'b000101;
 17'b00000110010110000 : data_comb = 6'b000110;
 17'b00000110010110001 : data_comb = 6'b000110;
 17'b00000110010110010 : data_comb = 6'b000110;
 17'b00000110010110011 : data_comb = 6'b000110;
 17'b00000110010110100 : data_comb = 6'b000110;
 17'b00000110010110101 : data_comb = 6'b000110;
 17'b00000110010110110 : data_comb = 6'b000110;
 17'b00000110010110111 : data_comb = 6'b000110;
 17'b00000110010111000 : data_comb = 6'b000110;
 17'b00000110010111001 : data_comb = 6'b000110;
 17'b00000110010111010 : data_comb = 6'b000110;
 17'b00000110010111011 : data_comb = 6'b000101;
 17'b00000110010111100 : data_comb = 6'b000101;
 17'b00000110010111101 : data_comb = 6'b000110;
 17'b00000110010111110 : data_comb = 6'b000110;
 17'b00000110010111111 : data_comb = 6'b000110;
 17'b00000110011000000 : data_comb = 6'b011001;
 17'b00000110011000001 : data_comb = 6'b111000;
 17'b00000110011000010 : data_comb = 6'b111000;
 17'b00000110011000011 : data_comb = 6'b000101;
 17'b00000110011000100 : data_comb = 6'b000110;
 17'b00000110011000101 : data_comb = 6'b000110;
 17'b00000110011000110 : data_comb = 6'b000110;
 17'b00000110011000111 : data_comb = 6'b101000;
 17'b00000110011001000 : data_comb = 6'b111000;
 17'b00000110011001001 : data_comb = 6'b111000;
 17'b00000110011001010 : data_comb = 6'b111000;
 17'b00000110011001011 : data_comb = 6'b111000;
 17'b00000110011001100 : data_comb = 6'b111000;
 17'b00000110011001101 : data_comb = 6'b111000;
 17'b00000110011001110 : data_comb = 6'b101000;
 17'b00000110011001111 : data_comb = 6'b101001;
 17'b00000110011010000 : data_comb = 6'b111000;
 17'b00000110011010001 : data_comb = 6'b111000;
 17'b00000110011010010 : data_comb = 6'b111000;
 17'b00000110011010011 : data_comb = 6'b111000;
 17'b00000110011010100 : data_comb = 6'b111000;
 17'b00000110011010101 : data_comb = 6'b111000;
 17'b00000110011010110 : data_comb = 6'b111000;
 17'b00000110011010111 : data_comb = 6'b111000;
 17'b00000110011011000 : data_comb = 6'b101001;
 17'b00000110011011001 : data_comb = 6'b000110;
 17'b00000110011011010 : data_comb = 6'b000110;
 17'b00000110011011011 : data_comb = 6'b000110;
 17'b00000110011011100 : data_comb = 6'b000110;
 17'b00000110011011101 : data_comb = 6'b000110;
 17'b00000110011011110 : data_comb = 6'b000110;
 17'b00000110011011111 : data_comb = 6'b000110;
 17'b00000110011100000 : data_comb = 6'b000101;
 17'b00000110011100001 : data_comb = 6'b000101;
 17'b00000110011100010 : data_comb = 6'b000101;
 17'b00000110011100011 : data_comb = 6'b000101;
 17'b00000110011100100 : data_comb = 6'b000110;
 17'b00000110011100101 : data_comb = 6'b000110;
 17'b00000110011100110 : data_comb = 6'b000110;
 17'b00000110011100111 : data_comb = 6'b000110;
 17'b00000110011101000 : data_comb = 6'b000101;
 17'b00000110011101001 : data_comb = 6'b000101;
 17'b00000110011101010 : data_comb = 6'b000101;
 17'b00000110011101011 : data_comb = 6'b000101;
 17'b00000110011101100 : data_comb = 6'b000101;
 17'b00000110011101101 : data_comb = 6'b000110;
 17'b00000110011101110 : data_comb = 6'b000110;
 17'b00000110011101111 : data_comb = 6'b000110;
 17'b00000110011110000 : data_comb = 6'b000110;
 17'b00000110011110001 : data_comb = 6'b000110;
 17'b00000110011110010 : data_comb = 6'b000110;
 17'b00000110011110011 : data_comb = 6'b000101;
 17'b00000110011110100 : data_comb = 6'b000101;
 17'b00000110011110101 : data_comb = 6'b000101;
 17'b00000110011110110 : data_comb = 6'b000101;
 17'b00000110011110111 : data_comb = 6'b000101;
 17'b00000110011111000 : data_comb = 6'b000101;
 17'b00000110011111001 : data_comb = 6'b000101;
 17'b00000110011111010 : data_comb = 6'b000110;
 17'b00000110011111011 : data_comb = 6'b000110;
 17'b00000110011111100 : data_comb = 6'b000110;
 17'b00000110011111101 : data_comb = 6'b000101;
 17'b00000110011111110 : data_comb = 6'b000101;
 17'b00000110011111111 : data_comb = 6'b000101;
 17'b00000110100000000 : data_comb = 6'b000101;
 17'b00000110100000001 : data_comb = 6'b000101;
 17'b00000110100000010 : data_comb = 6'b000110;
 17'b00000110100000011 : data_comb = 6'b000110;
 17'b00000110100000100 : data_comb = 6'b000110;
 17'b00000110100000101 : data_comb = 6'b000110;
 17'b00000110100000110 : data_comb = 6'b000110;
 17'b00000110100000111 : data_comb = 6'b000110;
 17'b00000110100001000 : data_comb = 6'b000110;
 17'b00000110100001001 : data_comb = 6'b000101;
 17'b00000110100001010 : data_comb = 6'b000101;
 17'b00000110100001011 : data_comb = 6'b000101;
 17'b00000110100001100 : data_comb = 6'b000101;
 17'b00000110100001101 : data_comb = 6'b000101;
 17'b00000110100001110 : data_comb = 6'b000101;
 17'b00000110100001111 : data_comb = 6'b011001;
 17'b00000110100010000 : data_comb = 6'b111000;
 17'b00000110100010001 : data_comb = 6'b111000;
 17'b00000110100010010 : data_comb = 6'b111000;
 17'b00000110100010011 : data_comb = 6'b111000;
 17'b00000110100010100 : data_comb = 6'b000101;
 17'b00000110100010101 : data_comb = 6'b000110;
 17'b00000110100010110 : data_comb = 6'b000110;
 17'b00000110100010111 : data_comb = 6'b000101;
 17'b00000110100011000 : data_comb = 6'b101000;
 17'b00000110100011001 : data_comb = 6'b111000;
 17'b00000110100011010 : data_comb = 6'b111000;
 17'b00000110100011011 : data_comb = 6'b111000;
 17'b00000110100011100 : data_comb = 6'b111000;
 17'b00000110100011101 : data_comb = 6'b111000;
 17'b00000110100011110 : data_comb = 6'b111000;
 17'b00000110100011111 : data_comb = 6'b111000;
 17'b00000110100100000 : data_comb = 6'b111000;
 17'b00000110100100001 : data_comb = 6'b111000;
 17'b00000110100100010 : data_comb = 6'b111000;
 17'b00000110100100011 : data_comb = 6'b111000;
 17'b00000110100100100 : data_comb = 6'b111000;
 17'b00000110100100101 : data_comb = 6'b111000;
 17'b00000110100100110 : data_comb = 6'b111000;
 17'b00000110100100111 : data_comb = 6'b111000;
 17'b00000110100101000 : data_comb = 6'b010101;
 17'b00000110100101001 : data_comb = 6'b000101;
 17'b00000110100101010 : data_comb = 6'b000110;
 17'b00000110100101011 : data_comb = 6'b000110;
 17'b00000110100101100 : data_comb = 6'b000110;
 17'b00000110100101101 : data_comb = 6'b000101;
 17'b00000110100101110 : data_comb = 6'b000101;
 17'b00000110100101111 : data_comb = 6'b000101;
 17'b00000110100110000 : data_comb = 6'b000101;
 17'b00000110100110001 : data_comb = 6'b000101;
 17'b00000110100110010 : data_comb = 6'b000101;
 17'b00000110100110011 : data_comb = 6'b000101;
 17'b00000110100110100 : data_comb = 6'b000101;
 17'b00000110100110101 : data_comb = 6'b000101;
 17'b00000110100110110 : data_comb = 6'b000110;
 17'b00000110100110111 : data_comb = 6'b000101;
 17'b00000110100111000 : data_comb = 6'b000101;
 17'b00000110100111001 : data_comb = 6'b000101;
 17'b00000110100111010 : data_comb = 6'b000101;
 17'b00000110100111011 : data_comb = 6'b000101;
 17'b00000110100111100 : data_comb = 6'b000101;
 17'b00000110100111101 : data_comb = 6'b000101;
 17'b00000110100111110 : data_comb = 6'b000110;
 17'b00000110100111111 : data_comb = 6'b000101;
 17'b00000110101000000 : data_comb = 6'b000101;
 17'b00000110101000001 : data_comb = 6'b000110;
 17'b00000110101000010 : data_comb = 6'b000110;
 17'b00000110101000011 : data_comb = 6'b000101;
 17'b00000110101000100 : data_comb = 6'b000101;
 17'b00000110101000101 : data_comb = 6'b000101;
 17'b00000110101000110 : data_comb = 6'b000101;
 17'b00000110101000111 : data_comb = 6'b000101;
 17'b00000110101001000 : data_comb = 6'b000101;
 17'b00000110101001001 : data_comb = 6'b000101;
 17'b00000110101001010 : data_comb = 6'b000101;
 17'b00000110101001011 : data_comb = 6'b000110;
 17'b00000110101001100 : data_comb = 6'b000101;
 17'b00000110101001101 : data_comb = 6'b000101;
 17'b00000110101001110 : data_comb = 6'b000101;
 17'b00000110101001111 : data_comb = 6'b000101;
 17'b00000110101010000 : data_comb = 6'b000101;
 17'b00000110101010001 : data_comb = 6'b000101;
 17'b00000110101010010 : data_comb = 6'b000101;
 17'b00000110101010011 : data_comb = 6'b000110;
 17'b00000110101010100 : data_comb = 6'b000101;
 17'b00000110101010101 : data_comb = 6'b000101;
 17'b00000110101010110 : data_comb = 6'b000101;
 17'b00000110101010111 : data_comb = 6'b000101;
 17'b00000110101011000 : data_comb = 6'b000101;
 17'b00000110101011001 : data_comb = 6'b000101;
 17'b00000110101011010 : data_comb = 6'b000101;
 17'b00000110101011011 : data_comb = 6'b000101;
 17'b00000110101011100 : data_comb = 6'b000101;
 17'b00000110101011101 : data_comb = 6'b000101;
 17'b00000110101011110 : data_comb = 6'b000101;
 17'b00000110101011111 : data_comb = 6'b011000;
 17'b00000110101100000 : data_comb = 6'b101000;
 17'b00000110101100001 : data_comb = 6'b111000;
 17'b00000110101100010 : data_comb = 6'b111000;
 17'b00000110101100011 : data_comb = 6'b111000;
 17'b00000110101100100 : data_comb = 6'b111000;
 17'b00000110101100101 : data_comb = 6'b011001;
 17'b00000110101100110 : data_comb = 6'b101000;
 17'b00000110101100111 : data_comb = 6'b111000;
 17'b00000110101101000 : data_comb = 6'b111000;
 17'b00000110101101001 : data_comb = 6'b111000;
 17'b00000110101101010 : data_comb = 6'b111000;
 17'b00000110101101011 : data_comb = 6'b111000;
 17'b00000110101101100 : data_comb = 6'b111000;
 17'b00000110101101101 : data_comb = 6'b111000;
 17'b00000110101101110 : data_comb = 6'b111000;
 17'b00000110101101111 : data_comb = 6'b111000;
 17'b00000110101110000 : data_comb = 6'b011001;
 17'b00000110101110001 : data_comb = 6'b111000;
 17'b00000110101110010 : data_comb = 6'b111000;
 17'b00000110101110011 : data_comb = 6'b111000;
 17'b00000110101110100 : data_comb = 6'b111000;
 17'b00000110101110101 : data_comb = 6'b111000;
 17'b00000110101110110 : data_comb = 6'b111000;
 17'b00000110101110111 : data_comb = 6'b111000;
 17'b00000110101111000 : data_comb = 6'b111000;
 17'b00000110101111001 : data_comb = 6'b011001;
 17'b00000110101111010 : data_comb = 6'b000110;
 17'b00000110101111011 : data_comb = 6'b000110;
 17'b00000110101111100 : data_comb = 6'b000101;
 17'b00000110101111101 : data_comb = 6'b000101;
 17'b00000110101111110 : data_comb = 6'b000101;
 17'b00000110101111111 : data_comb = 6'b000101;
 17'b00000110110000000 : data_comb = 6'b000101;
 17'b00000110110000001 : data_comb = 6'b000101;
 17'b00000110110000010 : data_comb = 6'b000101;
 17'b00000110110000011 : data_comb = 6'b000101;
 17'b00000110110000100 : data_comb = 6'b000101;
 17'b00000110110000101 : data_comb = 6'b000101;
 17'b00000110110000110 : data_comb = 6'b000101;
 17'b00000110110000111 : data_comb = 6'b000101;
 17'b00000110110001000 : data_comb = 6'b000101;
 17'b00000110110001001 : data_comb = 6'b000101;
 17'b00000110110001010 : data_comb = 6'b000101;
 17'b00000110110001011 : data_comb = 6'b000101;
 17'b00000110110001100 : data_comb = 6'b000101;
 17'b00000110110001101 : data_comb = 6'b000101;
 17'b00000110110001110 : data_comb = 6'b000101;
 17'b00000110110001111 : data_comb = 6'b000101;
 17'b00000110110010000 : data_comb = 6'b000101;
 17'b00000110110010001 : data_comb = 6'b000101;
 17'b00000110110010010 : data_comb = 6'b000110;
 17'b00000110110010011 : data_comb = 6'b000101;
 17'b00000110110010100 : data_comb = 6'b000101;
 17'b00000110110010101 : data_comb = 6'b000101;
 17'b00000110110010110 : data_comb = 6'b000101;
 17'b00000110110010111 : data_comb = 6'b000101;
 17'b00000110110011000 : data_comb = 6'b000101;
 17'b00000110110011001 : data_comb = 6'b000101;
 17'b00000110110011010 : data_comb = 6'b000101;
 17'b00000110110011011 : data_comb = 6'b000101;
 17'b00000110110011100 : data_comb = 6'b000101;
 17'b00000110110011101 : data_comb = 6'b000101;
 17'b00000110110011110 : data_comb = 6'b000101;
 17'b00000110110011111 : data_comb = 6'b000101;
 17'b00000110110100000 : data_comb = 6'b000101;
 17'b00000110110100001 : data_comb = 6'b000101;
 17'b00000110110100010 : data_comb = 6'b000101;
 17'b00000110110100011 : data_comb = 6'b000101;
 17'b00000110110100100 : data_comb = 6'b000101;
 17'b00000110110100101 : data_comb = 6'b000101;
 17'b00000110110100110 : data_comb = 6'b000101;
 17'b00000110110100111 : data_comb = 6'b000101;
 17'b00000110110101000 : data_comb = 6'b000101;
 17'b00000110110101001 : data_comb = 6'b000101;
 17'b00000110110101010 : data_comb = 6'b000101;
 17'b00000110110101011 : data_comb = 6'b000101;
 17'b00000110110101100 : data_comb = 6'b000101;
 17'b00000110110101101 : data_comb = 6'b000101;
 17'b00000110110101110 : data_comb = 6'b000101;
 17'b00000110110101111 : data_comb = 6'b000101;
 17'b00000110110110000 : data_comb = 6'b000101;
 17'b00000110110110001 : data_comb = 6'b010100;
 17'b00000110110110010 : data_comb = 6'b101000;
 17'b00000110110110011 : data_comb = 6'b111000;
 17'b00000110110110100 : data_comb = 6'b111000;
 17'b00000110110110101 : data_comb = 6'b111000;
 17'b00000110110110110 : data_comb = 6'b111000;
 17'b00000110110110111 : data_comb = 6'b111000;
 17'b00000110110111000 : data_comb = 6'b111000;
 17'b00000110110111001 : data_comb = 6'b111000;
 17'b00000110110111010 : data_comb = 6'b111000;
 17'b00000110110111011 : data_comb = 6'b111000;
 17'b00000110110111100 : data_comb = 6'b111000;
 17'b00000110110111101 : data_comb = 6'b101000;
 17'b00000110110111110 : data_comb = 6'b101000;
 17'b00000110110111111 : data_comb = 6'b101000;
 17'b00000110111000000 : data_comb = 6'b000110;
 17'b00000110111000001 : data_comb = 6'b000101;
 17'b00000110111000010 : data_comb = 6'b000101;
 17'b00000110111000011 : data_comb = 6'b101000;
 17'b00000110111000100 : data_comb = 6'b111000;
 17'b00000110111000101 : data_comb = 6'b111000;
 17'b00000110111000110 : data_comb = 6'b111000;
 17'b00000110111000111 : data_comb = 6'b111000;
 17'b00000110111001000 : data_comb = 6'b111000;
 17'b00000110111001001 : data_comb = 6'b111000;
 17'b00000110111001010 : data_comb = 6'b000101;
 17'b00000110111001011 : data_comb = 6'b000101;
 17'b00000110111001100 : data_comb = 6'b000101;
 17'b00000110111001101 : data_comb = 6'b000101;
 17'b00000110111001110 : data_comb = 6'b000101;
 17'b00000110111001111 : data_comb = 6'b000101;
 17'b00000110111010000 : data_comb = 6'b000101;
 17'b00000110111010001 : data_comb = 6'b000101;
 17'b00000110111010010 : data_comb = 6'b000101;
 17'b00000110111010011 : data_comb = 6'b000101;
 17'b00000110111010100 : data_comb = 6'b000101;
 17'b00000110111010101 : data_comb = 6'b000101;
 17'b00000110111010110 : data_comb = 6'b000101;
 17'b00000110111010111 : data_comb = 6'b000101;
 17'b00000110111011000 : data_comb = 6'b000101;
 17'b00000110111011001 : data_comb = 6'b000101;
 17'b00000110111011010 : data_comb = 6'b000101;
 17'b00000110111011011 : data_comb = 6'b000101;
 17'b00000110111011100 : data_comb = 6'b000101;
 17'b00000110111011101 : data_comb = 6'b000101;
 17'b00000110111011110 : data_comb = 6'b000101;
 17'b00000110111011111 : data_comb = 6'b000101;
 17'b00000110111100000 : data_comb = 6'b000101;
 17'b00000110111100001 : data_comb = 6'b000101;
 17'b00000110111100010 : data_comb = 6'b000101;
 17'b00000110111100011 : data_comb = 6'b000101;
 17'b00000110111100100 : data_comb = 6'b000101;
 17'b00000110111100101 : data_comb = 6'b000101;
 17'b00000110111100110 : data_comb = 6'b000101;
 17'b00000110111100111 : data_comb = 6'b000101;
 17'b00000110111101000 : data_comb = 6'b000101;
 17'b00000110111101001 : data_comb = 6'b000101;
 17'b00000110111101010 : data_comb = 6'b000101;
 17'b00000110111101011 : data_comb = 6'b000101;
 17'b00000110111101100 : data_comb = 6'b000101;
 17'b00000110111101101 : data_comb = 6'b000101;
 17'b00000110111101110 : data_comb = 6'b000101;
 17'b00000110111101111 : data_comb = 6'b000101;
 17'b00000110111110000 : data_comb = 6'b000101;
 17'b00000110111110001 : data_comb = 6'b000101;
 17'b00000110111110010 : data_comb = 6'b000101;
 17'b00000110111110011 : data_comb = 6'b000101;
 17'b00000110111110100 : data_comb = 6'b000101;
 17'b00000110111110101 : data_comb = 6'b000101;
 17'b00000110111110110 : data_comb = 6'b000101;
 17'b00000110111110111 : data_comb = 6'b000101;
 17'b00000110111111000 : data_comb = 6'b000101;
 17'b00000110111111001 : data_comb = 6'b000101;
 17'b00000110111111010 : data_comb = 6'b000101;
 17'b00000110111111011 : data_comb = 6'b000101;
 17'b00000110111111100 : data_comb = 6'b000101;
 17'b00000110111111101 : data_comb = 6'b000101;
 17'b00000110111111110 : data_comb = 6'b000101;
 17'b00000110111111111 : data_comb = 6'b000101;
 17'b00000111000000000 : data_comb = 6'b000101;
 17'b00000111000000001 : data_comb = 6'b000101;
 17'b00000111000000010 : data_comb = 6'b000101;
 17'b00000111000000011 : data_comb = 6'b010100;
 17'b00000111000000100 : data_comb = 6'b101000;
 17'b00000111000000101 : data_comb = 6'b111000;
 17'b00000111000000110 : data_comb = 6'b111000;
 17'b00000111000000111 : data_comb = 6'b111000;
 17'b00000111000001000 : data_comb = 6'b111000;
 17'b00000111000001001 : data_comb = 6'b111000;
 17'b00000111000001010 : data_comb = 6'b111000;
 17'b00000111000001011 : data_comb = 6'b111000;
 17'b00000111000001100 : data_comb = 6'b000101;
 17'b00000111000001101 : data_comb = 6'b000110;
 17'b00000111000001110 : data_comb = 6'b000110;
 17'b00000111000001111 : data_comb = 6'b000110;
 17'b00000111000010000 : data_comb = 6'b000110;
 17'b00000111000010001 : data_comb = 6'b000110;
 17'b00000111000010010 : data_comb = 6'b000110;
 17'b00000111000010011 : data_comb = 6'b000101;
 17'b00000111000010100 : data_comb = 6'b010101;
 17'b00000111000010101 : data_comb = 6'b010101;
 17'b00000111000010110 : data_comb = 6'b010101;
 17'b00000111000010111 : data_comb = 6'b010101;
 17'b00000111000011000 : data_comb = 6'b010101;
 17'b00000111000011001 : data_comb = 6'b010101;
 17'b00000111000011010 : data_comb = 6'b000101;
 17'b00000111000011011 : data_comb = 6'b000101;
 17'b00000111000011100 : data_comb = 6'b000101;
 17'b00000111000011101 : data_comb = 6'b000101;
 17'b00000111000011110 : data_comb = 6'b000101;
 17'b00000111000011111 : data_comb = 6'b000101;
 17'b00000111000100000 : data_comb = 6'b000101;
 17'b00000111000100001 : data_comb = 6'b000101;
 17'b00000111000100010 : data_comb = 6'b000101;
 17'b00000111000100011 : data_comb = 6'b000101;
 17'b00000111000100100 : data_comb = 6'b000101;
 17'b00000111000100101 : data_comb = 6'b000101;
 17'b00000111000100110 : data_comb = 6'b000101;
 17'b00000111000100111 : data_comb = 6'b000101;
 17'b00000111000101000 : data_comb = 6'b000101;
 17'b00000111000101001 : data_comb = 6'b000101;
 17'b00000111000101010 : data_comb = 6'b000101;
 17'b00000111000101011 : data_comb = 6'b000101;
 17'b00000111000101100 : data_comb = 6'b000101;
 17'b00000111000101101 : data_comb = 6'b000101;
 17'b00000111000101110 : data_comb = 6'b000101;
 17'b00000111000101111 : data_comb = 6'b000101;
 17'b00000111000110000 : data_comb = 6'b000101;
 17'b00000111000110001 : data_comb = 6'b000101;
 17'b00000111000110010 : data_comb = 6'b000101;
 17'b00000111000110011 : data_comb = 6'b000101;
 17'b00000111000110100 : data_comb = 6'b000101;
 17'b00000111000110101 : data_comb = 6'b000101;
 17'b00000111000110110 : data_comb = 6'b000101;
 17'b00000111000110111 : data_comb = 6'b000101;
 17'b00000111000111000 : data_comb = 6'b000101;
 17'b00000111000111001 : data_comb = 6'b000101;
 17'b00000111000111010 : data_comb = 6'b000101;
 17'b00000111000111011 : data_comb = 6'b000101;
 17'b00000111000111100 : data_comb = 6'b000101;
 17'b00000111000111101 : data_comb = 6'b000101;
 17'b00000111000111110 : data_comb = 6'b000101;
 17'b00000111000111111 : data_comb = 6'b000101;
 17'b00000111001000000 : data_comb = 6'b000101;
 17'b00000111001000001 : data_comb = 6'b000101;
 17'b00000111001000010 : data_comb = 6'b000101;
 17'b00000111001000011 : data_comb = 6'b000101;
 17'b00000111001000100 : data_comb = 6'b000101;
 17'b00000111001000101 : data_comb = 6'b000101;
 17'b00000111001000110 : data_comb = 6'b000101;
 17'b00000111001000111 : data_comb = 6'b000101;
 17'b00000111001001000 : data_comb = 6'b000101;
 17'b00000111001001001 : data_comb = 6'b000101;
 17'b00000111001001010 : data_comb = 6'b000101;
 17'b00000111001001011 : data_comb = 6'b000101;
 17'b00000111001001100 : data_comb = 6'b000101;
 17'b00000111001001101 : data_comb = 6'b000101;
 17'b00000111001001110 : data_comb = 6'b000101;
 17'b00000111001001111 : data_comb = 6'b000101;
 17'b00000111001010000 : data_comb = 6'b000101;
 17'b00000111001010001 : data_comb = 6'b000101;
 17'b00000111001010010 : data_comb = 6'b000101;
 17'b00000111001010011 : data_comb = 6'b000101;
 17'b00000111001010100 : data_comb = 6'b000101;
 17'b00000111001010101 : data_comb = 6'b000100;
 17'b00000111001010110 : data_comb = 6'b101000;
 17'b00000111001010111 : data_comb = 6'b000101;
 17'b00000111001011000 : data_comb = 6'b000110;
 17'b00000111001011001 : data_comb = 6'b000110;
 17'b00000111001011010 : data_comb = 6'b000110;
 17'b00000111001011011 : data_comb = 6'b000110;
 17'b00000111001011100 : data_comb = 6'b000110;
 17'b00000111001011101 : data_comb = 6'b000110;
 17'b00000111001011110 : data_comb = 6'b000110;
 17'b00000111001011111 : data_comb = 6'b000110;
 17'b00000111001100000 : data_comb = 6'b000110;
 17'b00000111001100001 : data_comb = 6'b000110;
 17'b00000111001100010 : data_comb = 6'b000110;
 17'b00000111001100011 : data_comb = 6'b000110;
 17'b00000111001100100 : data_comb = 6'b000110;
 17'b00000111001100101 : data_comb = 6'b000110;
 17'b00000111001100110 : data_comb = 6'b000110;
 17'b00000111001100111 : data_comb = 6'b000110;
 17'b00000111001101000 : data_comb = 6'b000110;
 17'b00000111001101001 : data_comb = 6'b000101;
 17'b00000111001101010 : data_comb = 6'b000101;
 17'b00000111001101011 : data_comb = 6'b000101;
 17'b00000111001101100 : data_comb = 6'b000101;
 17'b00000111001101101 : data_comb = 6'b000100;
 17'b00000111001101110 : data_comb = 6'b101000;
 17'b00000111001101111 : data_comb = 6'b101000;
 17'b00000111001110000 : data_comb = 6'b101000;
 17'b00000111001110001 : data_comb = 6'b101000;
 17'b00000111001110010 : data_comb = 6'b101000;
 17'b00000111001110011 : data_comb = 6'b101000;
 17'b00000111001110100 : data_comb = 6'b101000;
 17'b00000111001110101 : data_comb = 6'b101000;
 17'b00000111001110110 : data_comb = 6'b101000;
 17'b00000111001110111 : data_comb = 6'b101000;
 17'b00000111001111000 : data_comb = 6'b101000;
 17'b00000111001111001 : data_comb = 6'b101000;
 17'b00000111001111010 : data_comb = 6'b101000;
 17'b00000111001111011 : data_comb = 6'b101000;
 17'b00000111001111100 : data_comb = 6'b101000;
 17'b00000111001111101 : data_comb = 6'b101000;
 17'b00000111001111110 : data_comb = 6'b101000;
 17'b00000111001111111 : data_comb = 6'b101000;
 17'b00000111010000000 : data_comb = 6'b101000;
 17'b00000111010000001 : data_comb = 6'b101000;
 17'b00000111010000010 : data_comb = 6'b101000;
 17'b00000111010000011 : data_comb = 6'b101000;
 17'b00000111010000100 : data_comb = 6'b101000;
 17'b00000111010000101 : data_comb = 6'b101000;
 17'b00000111010000110 : data_comb = 6'b101000;
 17'b00000111010000111 : data_comb = 6'b101000;
 17'b00000111010001000 : data_comb = 6'b101000;
 17'b00000111010001001 : data_comb = 6'b101000;
 17'b00000111010001010 : data_comb = 6'b101000;
 17'b00000111010001011 : data_comb = 6'b101000;
 17'b00000111010001100 : data_comb = 6'b101000;
 17'b00000111010001101 : data_comb = 6'b101000;
 17'b00000111010001110 : data_comb = 6'b101000;
 17'b00000111010001111 : data_comb = 6'b101000;
 17'b00000111010010000 : data_comb = 6'b101000;
 17'b00000111010010001 : data_comb = 6'b101000;
 17'b00000111010010010 : data_comb = 6'b101000;
 17'b00000111010010011 : data_comb = 6'b101000;
 17'b00000111010010100 : data_comb = 6'b101000;
 17'b00000111010010101 : data_comb = 6'b101000;
 17'b00000111010010110 : data_comb = 6'b101000;
 17'b00000111010010111 : data_comb = 6'b101000;
 17'b00000111010011000 : data_comb = 6'b101000;
 17'b00000111010011001 : data_comb = 6'b101000;
 17'b00000111010011010 : data_comb = 6'b101000;
 17'b00000111010011011 : data_comb = 6'b101000;
 17'b00000111010011100 : data_comb = 6'b101000;
 17'b00000111010011101 : data_comb = 6'b101000;
 17'b00000111010011110 : data_comb = 6'b101000;
 17'b00000111010011111 : data_comb = 6'b101000;
 17'b00000111010100000 : data_comb = 6'b101000;
 17'b00000111010100001 : data_comb = 6'b101000;
 17'b00000111010100010 : data_comb = 6'b000100;
 17'b00000111010100011 : data_comb = 6'b000101;
 17'b00000111010100100 : data_comb = 6'b000101;
 17'b00000111010100101 : data_comb = 6'b000101;
 17'b00000111010100110 : data_comb = 6'b000101;
 17'b00000111010100111 : data_comb = 6'b000110;
 17'b00000111010101000 : data_comb = 6'b000110;
 17'b00000111010101001 : data_comb = 6'b000110;
 17'b00000111010101010 : data_comb = 6'b000110;
 17'b00000111010101011 : data_comb = 6'b000110;
 17'b00000111010101100 : data_comb = 6'b000110;
 17'b00000111010101101 : data_comb = 6'b000110;
 17'b00000111010101110 : data_comb = 6'b000110;
 17'b00000111010101111 : data_comb = 6'b000110;
 17'b00000111010110000 : data_comb = 6'b000110;
 17'b00000111010110001 : data_comb = 6'b000110;
 17'b00000111010110010 : data_comb = 6'b000110;
 17'b00000111010110011 : data_comb = 6'b000110;
 17'b00000111010110100 : data_comb = 6'b000110;
 17'b00000111010110101 : data_comb = 6'b000110;
 17'b00000111010110110 : data_comb = 6'b000110;
 17'b00000111010110111 : data_comb = 6'b000110;
 17'b00000111010111000 : data_comb = 6'b000110;
 17'b00000111010111001 : data_comb = 6'b000101;
 17'b00000111010111010 : data_comb = 6'b000101;
 17'b00000111010111011 : data_comb = 6'b000101;
 17'b00000111010111100 : data_comb = 6'b000100;
 17'b00000111010111101 : data_comb = 6'b011000;
 17'b00000111010111110 : data_comb = 6'b101000;
 17'b00000111010111111 : data_comb = 6'b101000;
 17'b00000111011000000 : data_comb = 6'b101000;
 17'b00000111011000001 : data_comb = 6'b101000;
 17'b00000111011000010 : data_comb = 6'b101000;
 17'b00000111011000011 : data_comb = 6'b101000;
 17'b00000111011000100 : data_comb = 6'b101000;
 17'b00000111011000101 : data_comb = 6'b101000;
 17'b00000111011000110 : data_comb = 6'b101000;
 17'b00000111011000111 : data_comb = 6'b101000;
 17'b00000111011001000 : data_comb = 6'b101000;
 17'b00000111011001001 : data_comb = 6'b101000;
 17'b00000111011001010 : data_comb = 6'b101000;
 17'b00000111011001011 : data_comb = 6'b101000;
 17'b00000111011001100 : data_comb = 6'b101000;
 17'b00000111011001101 : data_comb = 6'b101000;
 17'b00000111011001110 : data_comb = 6'b101000;
 17'b00000111011001111 : data_comb = 6'b101000;
 17'b00000111011010000 : data_comb = 6'b101000;
 17'b00000111011010001 : data_comb = 6'b101000;
 17'b00000111011010010 : data_comb = 6'b101000;
 17'b00000111011010011 : data_comb = 6'b101000;
 17'b00000111011010100 : data_comb = 6'b101000;
 17'b00000111011010101 : data_comb = 6'b101000;
 17'b00000111011010110 : data_comb = 6'b101000;
 17'b00000111011010111 : data_comb = 6'b101000;
 17'b00000111011011000 : data_comb = 6'b101000;
 17'b00000111011011001 : data_comb = 6'b101000;
 17'b00000111011011010 : data_comb = 6'b101000;
 17'b00000111011011011 : data_comb = 6'b101000;
 17'b00000111011011100 : data_comb = 6'b101000;
 17'b00000111011011101 : data_comb = 6'b101000;
 17'b00000111011011110 : data_comb = 6'b101000;
 17'b00000111011011111 : data_comb = 6'b101000;
 17'b00000111011100000 : data_comb = 6'b101000;
 17'b00000111011100001 : data_comb = 6'b101000;
 17'b00000111011100010 : data_comb = 6'b101000;
 17'b00000111011100011 : data_comb = 6'b101000;
 17'b00000111011100100 : data_comb = 6'b101000;
 17'b00000111011100101 : data_comb = 6'b101000;
 17'b00000111011100110 : data_comb = 6'b101000;
 17'b00000111011100111 : data_comb = 6'b101000;
 17'b00000111011101000 : data_comb = 6'b101000;
 17'b00000111011101001 : data_comb = 6'b101000;
 17'b00000111011101010 : data_comb = 6'b101000;
 17'b00000111011101011 : data_comb = 6'b101000;
 17'b00000111011101100 : data_comb = 6'b101000;
 17'b00000111011101101 : data_comb = 6'b101000;
 17'b00000111011101110 : data_comb = 6'b101000;
 17'b00000111011101111 : data_comb = 6'b101000;
 17'b00000111011110000 : data_comb = 6'b101000;
 17'b00000111011110001 : data_comb = 6'b101000;
 17'b00000111011110010 : data_comb = 6'b011000;
 17'b00000111011110011 : data_comb = 6'b000100;
 17'b00000111011110100 : data_comb = 6'b000101;
 17'b00000111011110101 : data_comb = 6'b000101;
 17'b00000111011110110 : data_comb = 6'b000101;
 17'b00000111011110111 : data_comb = 6'b000101;
 17'b00000111011111000 : data_comb = 6'b000110;
 17'b00000111011111001 : data_comb = 6'b000110;
 17'b00000111011111010 : data_comb = 6'b000110;
 17'b00000111011111011 : data_comb = 6'b000110;
 17'b00000111011111100 : data_comb = 6'b000110;
 17'b00000111011111101 : data_comb = 6'b000110;
 17'b00000111011111110 : data_comb = 6'b000110;
 17'b00000111011111111 : data_comb = 6'b000110;
 17'b00000111100000000 : data_comb = 6'b000110;
 17'b00000111100000001 : data_comb = 6'b000110;
 17'b00000111100000010 : data_comb = 6'b000110;
 17'b00000111100000011 : data_comb = 6'b011001;
 17'b00000111100000100 : data_comb = 6'b101001;
 17'b00000111100000101 : data_comb = 6'b011001;
 17'b00000111100000110 : data_comb = 6'b000110;
 17'b00000111100000111 : data_comb = 6'b000110;
 17'b00000111100001000 : data_comb = 6'b000110;
 17'b00000111100001001 : data_comb = 6'b000101;
 17'b00000111100001010 : data_comb = 6'b000101;
 17'b00000111100001011 : data_comb = 6'b000101;
 17'b00000111100001100 : data_comb = 6'b000100;
 17'b00000111100001101 : data_comb = 6'b011000;
 17'b00000111100001110 : data_comb = 6'b011000;
 17'b00000111100001111 : data_comb = 6'b011000;
 17'b00000111100010000 : data_comb = 6'b011000;
 17'b00000111100010001 : data_comb = 6'b011000;
 17'b00000111100010010 : data_comb = 6'b011000;
 17'b00000111100010011 : data_comb = 6'b011000;
 17'b00000111100010100 : data_comb = 6'b011000;
 17'b00000111100010101 : data_comb = 6'b011000;
 17'b00000111100010110 : data_comb = 6'b011000;
 17'b00000111100010111 : data_comb = 6'b011000;
 17'b00000111100011000 : data_comb = 6'b011000;
 17'b00000111100011001 : data_comb = 6'b011000;
 17'b00000111100011010 : data_comb = 6'b011000;
 17'b00000111100011011 : data_comb = 6'b011000;
 17'b00000111100011100 : data_comb = 6'b011000;
 17'b00000111100011101 : data_comb = 6'b011000;
 17'b00000111100011110 : data_comb = 6'b011000;
 17'b00000111100011111 : data_comb = 6'b011000;
 17'b00000111100100000 : data_comb = 6'b011000;
 17'b00000111100100001 : data_comb = 6'b011000;
 17'b00000111100100010 : data_comb = 6'b011000;
 17'b00000111100100011 : data_comb = 6'b011000;
 17'b00000111100100100 : data_comb = 6'b011000;
 17'b00000111100100101 : data_comb = 6'b011000;
 17'b00000111100100110 : data_comb = 6'b011000;
 17'b00000111100100111 : data_comb = 6'b011000;
 17'b00000111100101000 : data_comb = 6'b011000;
 17'b00000111100101001 : data_comb = 6'b011000;
 17'b00000111100101010 : data_comb = 6'b011000;
 17'b00000111100101011 : data_comb = 6'b011000;
 17'b00000111100101100 : data_comb = 6'b011000;
 17'b00000111100101101 : data_comb = 6'b011000;
 17'b00000111100101110 : data_comb = 6'b011000;
 17'b00000111100101111 : data_comb = 6'b011000;
 17'b00000111100110000 : data_comb = 6'b011000;
 17'b00000111100110001 : data_comb = 6'b011000;
 17'b00000111100110010 : data_comb = 6'b011000;
 17'b00000111100110011 : data_comb = 6'b011000;
 17'b00000111100110100 : data_comb = 6'b011000;
 17'b00000111100110101 : data_comb = 6'b011000;
 17'b00000111100110110 : data_comb = 6'b011000;
 17'b00000111100110111 : data_comb = 6'b011000;
 17'b00000111100111000 : data_comb = 6'b011000;
 17'b00000111100111001 : data_comb = 6'b011000;
 17'b00000111100111010 : data_comb = 6'b011000;
 17'b00000111100111011 : data_comb = 6'b011000;
 17'b00000111100111100 : data_comb = 6'b011000;
 17'b00000111100111101 : data_comb = 6'b011000;
 17'b00000111100111110 : data_comb = 6'b011000;
 17'b00000111100111111 : data_comb = 6'b011000;
 17'b00000111101000000 : data_comb = 6'b011000;
 17'b00000111101000001 : data_comb = 6'b011000;
 17'b00000111101000010 : data_comb = 6'b011000;
 17'b00000111101000011 : data_comb = 6'b010100;
 17'b00000111101000100 : data_comb = 6'b000101;
 17'b00000111101000101 : data_comb = 6'b000101;
 17'b00000111101000110 : data_comb = 6'b000101;
 17'b00000111101000111 : data_comb = 6'b000101;
 17'b00000111101001000 : data_comb = 6'b000110;
 17'b00000111101001001 : data_comb = 6'b000110;
 17'b00000111101001010 : data_comb = 6'b000101;
 17'b00000111101001011 : data_comb = 6'b011001;
 17'b00000111101001100 : data_comb = 6'b011001;
 17'b00000111101001101 : data_comb = 6'b000101;
 17'b00000111101001110 : data_comb = 6'b000110;
 17'b00000111101001111 : data_comb = 6'b000110;
 17'b00000111101010000 : data_comb = 6'b000110;
 17'b00000111101010001 : data_comb = 6'b000110;
 17'b00000111101010010 : data_comb = 6'b011001;
 17'b00000111101010011 : data_comb = 6'b111000;
 17'b00000111101010100 : data_comb = 6'b111000;
 17'b00000111101010101 : data_comb = 6'b111000;
 17'b00000111101010110 : data_comb = 6'b011001;
 17'b00000111101010111 : data_comb = 6'b000110;
 17'b00000111101011000 : data_comb = 6'b000101;
 17'b00000111101011001 : data_comb = 6'b000101;
 17'b00000111101011010 : data_comb = 6'b000101;
 17'b00000111101011011 : data_comb = 6'b000101;
 17'b00000111101011100 : data_comb = 6'b000100;
 17'b00000111101011101 : data_comb = 6'b011000;
 17'b00000111101011110 : data_comb = 6'b011000;
 17'b00000111101011111 : data_comb = 6'b011000;
 17'b00000111101100000 : data_comb = 6'b011000;
 17'b00000111101100001 : data_comb = 6'b011000;
 17'b00000111101100010 : data_comb = 6'b011000;
 17'b00000111101100011 : data_comb = 6'b011000;
 17'b00000111101100100 : data_comb = 6'b011000;
 17'b00000111101100101 : data_comb = 6'b011000;
 17'b00000111101100110 : data_comb = 6'b011000;
 17'b00000111101100111 : data_comb = 6'b011000;
 17'b00000111101101000 : data_comb = 6'b011000;
 17'b00000111101101001 : data_comb = 6'b011000;
 17'b00000111101101010 : data_comb = 6'b011000;
 17'b00000111101101011 : data_comb = 6'b011000;
 17'b00000111101101100 : data_comb = 6'b011000;
 17'b00000111101101101 : data_comb = 6'b011000;
 17'b00000111101101110 : data_comb = 6'b011000;
 17'b00000111101101111 : data_comb = 6'b011000;
 17'b00000111101110000 : data_comb = 6'b011000;
 17'b00000111101110001 : data_comb = 6'b011000;
 17'b00000111101110010 : data_comb = 6'b011000;
 17'b00000111101110011 : data_comb = 6'b011000;
 17'b00000111101110100 : data_comb = 6'b011000;
 17'b00000111101110101 : data_comb = 6'b011000;
 17'b00000111101110110 : data_comb = 6'b011000;
 17'b00000111101110111 : data_comb = 6'b011000;
 17'b00000111101111000 : data_comb = 6'b011000;
 17'b00000111101111001 : data_comb = 6'b011000;
 17'b00000111101111010 : data_comb = 6'b011000;
 17'b00000111101111011 : data_comb = 6'b011000;
 17'b00000111101111100 : data_comb = 6'b011000;
 17'b00000111101111101 : data_comb = 6'b011000;
 17'b00000111101111110 : data_comb = 6'b011000;
 17'b00000111101111111 : data_comb = 6'b011000;
 17'b00000111110000000 : data_comb = 6'b011000;
 17'b00000111110000001 : data_comb = 6'b011000;
 17'b00000111110000010 : data_comb = 6'b011000;
 17'b00000111110000011 : data_comb = 6'b011000;
 17'b00000111110000100 : data_comb = 6'b011000;
 17'b00000111110000101 : data_comb = 6'b011000;
 17'b00000111110000110 : data_comb = 6'b011000;
 17'b00000111110000111 : data_comb = 6'b011000;
 17'b00000111110001000 : data_comb = 6'b011000;
 17'b00000111110001001 : data_comb = 6'b011000;
 17'b00000111110001010 : data_comb = 6'b011000;
 17'b00000111110001011 : data_comb = 6'b011000;
 17'b00000111110001100 : data_comb = 6'b011000;
 17'b00000111110001101 : data_comb = 6'b011000;
 17'b00000111110001110 : data_comb = 6'b011000;
 17'b00000111110001111 : data_comb = 6'b011000;
 17'b00000111110010000 : data_comb = 6'b011000;
 17'b00000111110010001 : data_comb = 6'b011000;
 17'b00000111110010010 : data_comb = 6'b011000;
 17'b00000111110010011 : data_comb = 6'b000100;
 17'b00000111110010100 : data_comb = 6'b000101;
 17'b00000111110010101 : data_comb = 6'b000101;
 17'b00000111110010110 : data_comb = 6'b000101;
 17'b00000111110010111 : data_comb = 6'b000101;
 17'b00000111110011000 : data_comb = 6'b000110;
 17'b00000111110011001 : data_comb = 6'b000101;
 17'b00000111110011010 : data_comb = 6'b101000;
 17'b00000111110011011 : data_comb = 6'b111000;
 17'b00000111110011100 : data_comb = 6'b111000;
 17'b00000111110011101 : data_comb = 6'b101000;
 17'b00000111110011110 : data_comb = 6'b000101;
 17'b00000111110011111 : data_comb = 6'b000110;
 17'b00000111110100000 : data_comb = 6'b011001;
 17'b00000111110100001 : data_comb = 6'b101001;
 17'b00000111110100010 : data_comb = 6'b111000;
 17'b00000111110100011 : data_comb = 6'b111000;
 17'b00000111110100100 : data_comb = 6'b111000;
 17'b00000111110100101 : data_comb = 6'b111000;
 17'b00000111110100110 : data_comb = 6'b111000;
 17'b00000111110100111 : data_comb = 6'b000110;
 17'b00000111110101000 : data_comb = 6'b000101;
 17'b00000111110101001 : data_comb = 6'b000101;
 17'b00000111110101010 : data_comb = 6'b000101;
 17'b00000111110101011 : data_comb = 6'b000101;
 17'b00000111110101100 : data_comb = 6'b000100;
 17'b00000111110101101 : data_comb = 6'b011000;
 17'b00000111110101110 : data_comb = 6'b000100;
 17'b00000111110101111 : data_comb = 6'b000101;
 17'b00000111110110000 : data_comb = 6'b000100;
 17'b00000111110110001 : data_comb = 6'b011000;
 17'b00000111110110010 : data_comb = 6'b000100;
 17'b00000111110110011 : data_comb = 6'b000101;
 17'b00000111110110100 : data_comb = 6'b000100;
 17'b00000111110110101 : data_comb = 6'b011000;
 17'b00000111110110110 : data_comb = 6'b011000;
 17'b00000111110110111 : data_comb = 6'b000100;
 17'b00000111110111000 : data_comb = 6'b000101;
 17'b00000111110111001 : data_comb = 6'b000101;
 17'b00000111110111010 : data_comb = 6'b000100;
 17'b00000111110111011 : data_comb = 6'b011000;
 17'b00000111110111100 : data_comb = 6'b011000;
 17'b00000111110111101 : data_comb = 6'b011000;
 17'b00000111110111110 : data_comb = 6'b000100;
 17'b00000111110111111 : data_comb = 6'b000101;
 17'b00000111111000000 : data_comb = 6'b000101;
 17'b00000111111000001 : data_comb = 6'b000100;
 17'b00000111111000010 : data_comb = 6'b011000;
 17'b00000111111000011 : data_comb = 6'b011000;
 17'b00000111111000100 : data_comb = 6'b000100;
 17'b00000111111000101 : data_comb = 6'b000101;
 17'b00000111111000110 : data_comb = 6'b000100;
 17'b00000111111000111 : data_comb = 6'b011000;
 17'b00000111111001000 : data_comb = 6'b011000;
 17'b00000111111001001 : data_comb = 6'b000100;
 17'b00000111111001010 : data_comb = 6'b000101;
 17'b00000111111001011 : data_comb = 6'b000101;
 17'b00000111111001100 : data_comb = 6'b000101;
 17'b00000111111001101 : data_comb = 6'b011000;
 17'b00000111111001110 : data_comb = 6'b011000;
 17'b00000111111001111 : data_comb = 6'b011000;
 17'b00000111111010000 : data_comb = 6'b011000;
 17'b00000111111010001 : data_comb = 6'b000100;
 17'b00000111111010010 : data_comb = 6'b000101;
 17'b00000111111010011 : data_comb = 6'b000100;
 17'b00000111111010100 : data_comb = 6'b011000;
 17'b00000111111010101 : data_comb = 6'b011000;
 17'b00000111111010110 : data_comb = 6'b000100;
 17'b00000111111010111 : data_comb = 6'b000101;
 17'b00000111111011000 : data_comb = 6'b000100;
 17'b00000111111011001 : data_comb = 6'b011000;
 17'b00000111111011010 : data_comb = 6'b010100;
 17'b00000111111011011 : data_comb = 6'b000101;
 17'b00000111111011100 : data_comb = 6'b000101;
 17'b00000111111011101 : data_comb = 6'b000100;
 17'b00000111111011110 : data_comb = 6'b011000;
 17'b00000111111011111 : data_comb = 6'b000100;
 17'b00000111111100000 : data_comb = 6'b000101;
 17'b00000111111100001 : data_comb = 6'b000101;
 17'b00000111111100010 : data_comb = 6'b011000;
 17'b00000111111100011 : data_comb = 6'b000100;
 17'b00000111111100100 : data_comb = 6'b000101;
 17'b00000111111100101 : data_comb = 6'b000101;
 17'b00000111111100110 : data_comb = 6'b000101;
 17'b00000111111100111 : data_comb = 6'b000101;
 17'b00000111111101000 : data_comb = 6'b000101;
 17'b00000111111101001 : data_comb = 6'b111000;
 17'b00000111111101010 : data_comb = 6'b111000;
 17'b00000111111101011 : data_comb = 6'b111000;
 17'b00000111111101100 : data_comb = 6'b111000;
 17'b00000111111101101 : data_comb = 6'b111000;
 17'b00000111111101110 : data_comb = 6'b101000;
 17'b00000111111101111 : data_comb = 6'b000101;
 17'b00000111111110000 : data_comb = 6'b111000;
 17'b00000111111110001 : data_comb = 6'b111000;
 17'b00000111111110010 : data_comb = 6'b111000;
 17'b00000111111110011 : data_comb = 6'b111000;
 17'b00000111111110100 : data_comb = 6'b111000;
 17'b00000111111110101 : data_comb = 6'b111000;
 17'b00000111111110110 : data_comb = 6'b111000;
 17'b00000111111110111 : data_comb = 6'b000100;
 17'b00000111111111000 : data_comb = 6'b000101;
 17'b00000111111111001 : data_comb = 6'b000101;
 17'b00000111111111010 : data_comb = 6'b000101;
 17'b00000111111111011 : data_comb = 6'b000101;
 17'b00000111111111100 : data_comb = 6'b000000;
 17'b00000111111111101 : data_comb = 6'b000000;
 17'b00000111111111110 : data_comb = 6'b000000;
 17'b00000111111111111 : data_comb = 6'b000000;
 17'b00001000000000000 : data_comb = 6'b000000;
 17'b00001000000000001 : data_comb = 6'b000000;
 17'b00001000000000010 : data_comb = 6'b000000;
 17'b00001000000000011 : data_comb = 6'b000000;
 17'b00001000000000100 : data_comb = 6'b000000;
 17'b00001000000000101 : data_comb = 6'b000000;
 17'b00001000000000110 : data_comb = 6'b000000;
 17'b00001000000000111 : data_comb = 6'b000000;
 17'b00001000000001000 : data_comb = 6'b000000;
 17'b00001000000001001 : data_comb = 6'b000000;
 17'b00001000000001010 : data_comb = 6'b000000;
 17'b00001000000001011 : data_comb = 6'b000000;
 17'b00001000000001100 : data_comb = 6'b000000;
 17'b00001000000001101 : data_comb = 6'b000000;
 17'b00001000000001110 : data_comb = 6'b000000;
 17'b00001000000001111 : data_comb = 6'b000000;
 17'b00001000000010000 : data_comb = 6'b000000;
 17'b00001000000010001 : data_comb = 6'b000000;
 17'b00001000000010010 : data_comb = 6'b000000;
 17'b00001000000010011 : data_comb = 6'b000000;
 17'b00001000000010100 : data_comb = 6'b000000;
 17'b00001000000010101 : data_comb = 6'b000000;
 17'b00001000000010110 : data_comb = 6'b000000;
 17'b00001000000010111 : data_comb = 6'b000000;
 17'b00001000000011000 : data_comb = 6'b000000;
 17'b00001000000011001 : data_comb = 6'b000000;
 17'b00001000000011010 : data_comb = 6'b000000;
 17'b00001000000011011 : data_comb = 6'b000000;
 17'b00001000000011100 : data_comb = 6'b000000;
 17'b00001000000011101 : data_comb = 6'b000000;
 17'b00001000000011110 : data_comb = 6'b000000;
 17'b00001000000011111 : data_comb = 6'b000000;
 17'b00001000000100000 : data_comb = 6'b000000;
 17'b00001000000100001 : data_comb = 6'b000000;
 17'b00001000000100010 : data_comb = 6'b000000;
 17'b00001000000100011 : data_comb = 6'b000000;
 17'b00001000000100100 : data_comb = 6'b000000;
 17'b00001000000100101 : data_comb = 6'b000000;
 17'b00001000000100110 : data_comb = 6'b000000;
 17'b00001000000100111 : data_comb = 6'b000000;
 17'b00001000000101000 : data_comb = 6'b000000;
 17'b00001000000101001 : data_comb = 6'b000000;
 17'b00001000000101010 : data_comb = 6'b000000;
 17'b00001000000101011 : data_comb = 6'b000000;
 17'b00001000000101100 : data_comb = 6'b000000;
 17'b00001000000101101 : data_comb = 6'b000000;
 17'b00001000000101110 : data_comb = 6'b000000;
 17'b00001000000101111 : data_comb = 6'b000000;
 17'b00001000000110000 : data_comb = 6'b000000;
 17'b00001000000110001 : data_comb = 6'b000000;
 17'b00001000000110010 : data_comb = 6'b000000;
 17'b00001000000110011 : data_comb = 6'b000000;
 17'b00001000000110100 : data_comb = 6'b000101;
 17'b00001000000110101 : data_comb = 6'b000101;
 17'b00001000000110110 : data_comb = 6'b000101;
 17'b00001000000110111 : data_comb = 6'b000101;
 17'b00001000000111000 : data_comb = 6'b000101;
 17'b00001000000111001 : data_comb = 6'b111000;
 17'b00001000000111010 : data_comb = 6'b111000;
 17'b00001000000111011 : data_comb = 6'b111000;
 17'b00001000000111100 : data_comb = 6'b111000;
 17'b00001000000111101 : data_comb = 6'b111000;
 17'b00001000000111110 : data_comb = 6'b111000;
 17'b00001000000111111 : data_comb = 6'b111000;
 17'b00001000001000000 : data_comb = 6'b111000;
 17'b00001000001000001 : data_comb = 6'b111000;
 17'b00001000001000010 : data_comb = 6'b111000;
 17'b00001000001000011 : data_comb = 6'b111000;
 17'b00001000001000100 : data_comb = 6'b111000;
 17'b00001000001000101 : data_comb = 6'b111000;
 17'b00001000001000110 : data_comb = 6'b111000;
 17'b00001000001000111 : data_comb = 6'b010100;
 17'b00001000001001000 : data_comb = 6'b000101;
 17'b00001000001001001 : data_comb = 6'b000101;
 17'b00001000001001010 : data_comb = 6'b000101;
 17'b00001000001001011 : data_comb = 6'b000101;
 17'b00001000001001100 : data_comb = 6'b000001;
 17'b00001000001001101 : data_comb = 6'b000000;
 17'b00001000001001110 : data_comb = 6'b000000;
 17'b00001000001001111 : data_comb = 6'b000000;
 17'b00001000001010000 : data_comb = 6'b010000;
 17'b00001000001010001 : data_comb = 6'b010000;
 17'b00001000001010010 : data_comb = 6'b010000;
 17'b00001000001010011 : data_comb = 6'b010000;
 17'b00001000001010100 : data_comb = 6'b010000;
 17'b00001000001010101 : data_comb = 6'b000000;
 17'b00001000001010110 : data_comb = 6'b000000;
 17'b00001000001010111 : data_comb = 6'b000000;
 17'b00001000001011000 : data_comb = 6'b000000;
 17'b00001000001011001 : data_comb = 6'b000000;
 17'b00001000001011010 : data_comb = 6'b000000;
 17'b00001000001011011 : data_comb = 6'b000000;
 17'b00001000001011100 : data_comb = 6'b000000;
 17'b00001000001011101 : data_comb = 6'b000000;
 17'b00001000001011110 : data_comb = 6'b010000;
 17'b00001000001011111 : data_comb = 6'b010000;
 17'b00001000001100000 : data_comb = 6'b010000;
 17'b00001000001100001 : data_comb = 6'b000000;
 17'b00001000001100010 : data_comb = 6'b000000;
 17'b00001000001100011 : data_comb = 6'b010000;
 17'b00001000001100100 : data_comb = 6'b010000;
 17'b00001000001100101 : data_comb = 6'b010000;
 17'b00001000001100110 : data_comb = 6'b010000;
 17'b00001000001100111 : data_comb = 6'b010000;
 17'b00001000001101000 : data_comb = 6'b000000;
 17'b00001000001101001 : data_comb = 6'b000000;
 17'b00001000001101010 : data_comb = 6'b000000;
 17'b00001000001101011 : data_comb = 6'b000000;
 17'b00001000001101100 : data_comb = 6'b010000;
 17'b00001000001101101 : data_comb = 6'b010000;
 17'b00001000001101110 : data_comb = 6'b000000;
 17'b00001000001101111 : data_comb = 6'b000000;
 17'b00001000001110000 : data_comb = 6'b010000;
 17'b00001000001110001 : data_comb = 6'b010000;
 17'b00001000001110010 : data_comb = 6'b010000;
 17'b00001000001110011 : data_comb = 6'b000000;
 17'b00001000001110100 : data_comb = 6'b000000;
 17'b00001000001110101 : data_comb = 6'b000000;
 17'b00001000001110110 : data_comb = 6'b000000;
 17'b00001000001110111 : data_comb = 6'b010000;
 17'b00001000001111000 : data_comb = 6'b010000;
 17'b00001000001111001 : data_comb = 6'b010000;
 17'b00001000001111010 : data_comb = 6'b010000;
 17'b00001000001111011 : data_comb = 6'b000000;
 17'b00001000001111100 : data_comb = 6'b000000;
 17'b00001000001111101 : data_comb = 6'b010000;
 17'b00001000001111110 : data_comb = 6'b010000;
 17'b00001000001111111 : data_comb = 6'b010000;
 17'b00001000010000000 : data_comb = 6'b000000;
 17'b00001000010000001 : data_comb = 6'b000000;
 17'b00001000010000010 : data_comb = 6'b000000;
 17'b00001000010000011 : data_comb = 6'b000001;
 17'b00001000010000100 : data_comb = 6'b000101;
 17'b00001000010000101 : data_comb = 6'b000101;
 17'b00001000010000110 : data_comb = 6'b000101;
 17'b00001000010000111 : data_comb = 6'b000101;
 17'b00001000010001000 : data_comb = 6'b010100;
 17'b00001000010001001 : data_comb = 6'b111000;
 17'b00001000010001010 : data_comb = 6'b111000;
 17'b00001000010001011 : data_comb = 6'b111000;
 17'b00001000010001100 : data_comb = 6'b111000;
 17'b00001000010001101 : data_comb = 6'b111000;
 17'b00001000010001110 : data_comb = 6'b111000;
 17'b00001000010001111 : data_comb = 6'b111000;
 17'b00001000010010000 : data_comb = 6'b111000;
 17'b00001000010010001 : data_comb = 6'b101000;
 17'b00001000010010010 : data_comb = 6'b011000;
 17'b00001000010010011 : data_comb = 6'b000101;
 17'b00001000010010100 : data_comb = 6'b000101;
 17'b00001000010010101 : data_comb = 6'b011000;
 17'b00001000010010110 : data_comb = 6'b101000;
 17'b00001000010010111 : data_comb = 6'b111000;
 17'b00001000010011000 : data_comb = 6'b000101;
 17'b00001000010011001 : data_comb = 6'b000101;
 17'b00001000010011010 : data_comb = 6'b000101;
 17'b00001000010011011 : data_comb = 6'b000101;
 17'b00001000010011100 : data_comb = 6'b000001;
 17'b00001000010011101 : data_comb = 6'b000001;
 17'b00001000010011110 : data_comb = 6'b000000;
 17'b00001000010011111 : data_comb = 6'b000000;
 17'b00001000010100000 : data_comb = 6'b010000;
 17'b00001000010100001 : data_comb = 6'b010000;
 17'b00001000010100010 : data_comb = 6'b010000;
 17'b00001000010100011 : data_comb = 6'b010000;
 17'b00001000010100100 : data_comb = 6'b010000;
 17'b00001000010100101 : data_comb = 6'b000000;
 17'b00001000010100110 : data_comb = 6'b000000;
 17'b00001000010100111 : data_comb = 6'b010000;
 17'b00001000010101000 : data_comb = 6'b010000;
 17'b00001000010101001 : data_comb = 6'b010000;
 17'b00001000010101010 : data_comb = 6'b010000;
 17'b00001000010101011 : data_comb = 6'b010000;
 17'b00001000010101100 : data_comb = 6'b000000;
 17'b00001000010101101 : data_comb = 6'b000000;
 17'b00001000010101110 : data_comb = 6'b010000;
 17'b00001000010101111 : data_comb = 6'b010000;
 17'b00001000010110000 : data_comb = 6'b010000;
 17'b00001000010110001 : data_comb = 6'b000000;
 17'b00001000010110010 : data_comb = 6'b000000;
 17'b00001000010110011 : data_comb = 6'b010000;
 17'b00001000010110100 : data_comb = 6'b010000;
 17'b00001000010110101 : data_comb = 6'b010000;
 17'b00001000010110110 : data_comb = 6'b010000;
 17'b00001000010110111 : data_comb = 6'b010000;
 17'b00001000010111000 : data_comb = 6'b010000;
 17'b00001000010111001 : data_comb = 6'b000000;
 17'b00001000010111010 : data_comb = 6'b000000;
 17'b00001000010111011 : data_comb = 6'b010000;
 17'b00001000010111100 : data_comb = 6'b010000;
 17'b00001000010111101 : data_comb = 6'b010000;
 17'b00001000010111110 : data_comb = 6'b000000;
 17'b00001000010111111 : data_comb = 6'b000000;
 17'b00001000011000000 : data_comb = 6'b010000;
 17'b00001000011000001 : data_comb = 6'b010000;
 17'b00001000011000010 : data_comb = 6'b010000;
 17'b00001000011000011 : data_comb = 6'b010000;
 17'b00001000011000100 : data_comb = 6'b000000;
 17'b00001000011000101 : data_comb = 6'b000000;
 17'b00001000011000110 : data_comb = 6'b000000;
 17'b00001000011000111 : data_comb = 6'b010000;
 17'b00001000011001000 : data_comb = 6'b010000;
 17'b00001000011001001 : data_comb = 6'b010000;
 17'b00001000011001010 : data_comb = 6'b010000;
 17'b00001000011001011 : data_comb = 6'b000000;
 17'b00001000011001100 : data_comb = 6'b010000;
 17'b00001000011001101 : data_comb = 6'b010000;
 17'b00001000011001110 : data_comb = 6'b010000;
 17'b00001000011001111 : data_comb = 6'b010000;
 17'b00001000011010000 : data_comb = 6'b000000;
 17'b00001000011010001 : data_comb = 6'b000000;
 17'b00001000011010010 : data_comb = 6'b000000;
 17'b00001000011010011 : data_comb = 6'b000001;
 17'b00001000011010100 : data_comb = 6'b000101;
 17'b00001000011010101 : data_comb = 6'b000101;
 17'b00001000011010110 : data_comb = 6'b000101;
 17'b00001000011010111 : data_comb = 6'b000101;
 17'b00001000011011000 : data_comb = 6'b000101;
 17'b00001000011011001 : data_comb = 6'b111000;
 17'b00001000011011010 : data_comb = 6'b111000;
 17'b00001000011011011 : data_comb = 6'b111000;
 17'b00001000011011100 : data_comb = 6'b111000;
 17'b00001000011011101 : data_comb = 6'b101000;
 17'b00001000011011110 : data_comb = 6'b010101;
 17'b00001000011011111 : data_comb = 6'b101000;
 17'b00001000011100000 : data_comb = 6'b000101;
 17'b00001000011100001 : data_comb = 6'b000101;
 17'b00001000011100010 : data_comb = 6'b000101;
 17'b00001000011100011 : data_comb = 6'b000101;
 17'b00001000011100100 : data_comb = 6'b000101;
 17'b00001000011100101 : data_comb = 6'b000101;
 17'b00001000011100110 : data_comb = 6'b000101;
 17'b00001000011100111 : data_comb = 6'b101000;
 17'b00001000011101000 : data_comb = 6'b010100;
 17'b00001000011101001 : data_comb = 6'b000101;
 17'b00001000011101010 : data_comb = 6'b000001;
 17'b00001000011101011 : data_comb = 6'b000001;
 17'b00001000011101100 : data_comb = 6'b000001;
 17'b00001000011101101 : data_comb = 6'b000001;
 17'b00001000011101110 : data_comb = 6'b000000;
 17'b00001000011101111 : data_comb = 6'b000000;
 17'b00001000011110000 : data_comb = 6'b010000;
 17'b00001000011110001 : data_comb = 6'b010000;
 17'b00001000011110010 : data_comb = 6'b010000;
 17'b00001000011110011 : data_comb = 6'b010000;
 17'b00001000011110100 : data_comb = 6'b010000;
 17'b00001000011110101 : data_comb = 6'b000000;
 17'b00001000011110110 : data_comb = 6'b000000;
 17'b00001000011110111 : data_comb = 6'b010000;
 17'b00001000011111000 : data_comb = 6'b010000;
 17'b00001000011111001 : data_comb = 6'b010000;
 17'b00001000011111010 : data_comb = 6'b010000;
 17'b00001000011111011 : data_comb = 6'b010000;
 17'b00001000011111100 : data_comb = 6'b000000;
 17'b00001000011111101 : data_comb = 6'b000000;
 17'b00001000011111110 : data_comb = 6'b010000;
 17'b00001000011111111 : data_comb = 6'b010000;
 17'b00001000100000000 : data_comb = 6'b010000;
 17'b00001000100000001 : data_comb = 6'b000000;
 17'b00001000100000010 : data_comb = 6'b000000;
 17'b00001000100000011 : data_comb = 6'b010000;
 17'b00001000100000100 : data_comb = 6'b010000;
 17'b00001000100000101 : data_comb = 6'b010000;
 17'b00001000100000110 : data_comb = 6'b010000;
 17'b00001000100000111 : data_comb = 6'b010000;
 17'b00001000100001000 : data_comb = 6'b010000;
 17'b00001000100001001 : data_comb = 6'b010000;
 17'b00001000100001010 : data_comb = 6'b000000;
 17'b00001000100001011 : data_comb = 6'b010000;
 17'b00001000100001100 : data_comb = 6'b010000;
 17'b00001000100001101 : data_comb = 6'b010000;
 17'b00001000100001110 : data_comb = 6'b000000;
 17'b00001000100001111 : data_comb = 6'b000000;
 17'b00001000100010000 : data_comb = 6'b010000;
 17'b00001000100010001 : data_comb = 6'b010000;
 17'b00001000100010010 : data_comb = 6'b010000;
 17'b00001000100010011 : data_comb = 6'b010000;
 17'b00001000100010100 : data_comb = 6'b010000;
 17'b00001000100010101 : data_comb = 6'b010000;
 17'b00001000100010110 : data_comb = 6'b000000;
 17'b00001000100010111 : data_comb = 6'b010000;
 17'b00001000100011000 : data_comb = 6'b010000;
 17'b00001000100011001 : data_comb = 6'b010000;
 17'b00001000100011010 : data_comb = 6'b010000;
 17'b00001000100011011 : data_comb = 6'b000000;
 17'b00001000100011100 : data_comb = 6'b010000;
 17'b00001000100011101 : data_comb = 6'b010000;
 17'b00001000100011110 : data_comb = 6'b010000;
 17'b00001000100011111 : data_comb = 6'b010000;
 17'b00001000100100000 : data_comb = 6'b000000;
 17'b00001000100100001 : data_comb = 6'b000000;
 17'b00001000100100010 : data_comb = 6'b000001;
 17'b00001000100100011 : data_comb = 6'b000001;
 17'b00001000100100100 : data_comb = 6'b000001;
 17'b00001000100100101 : data_comb = 6'b000001;
 17'b00001000100100110 : data_comb = 6'b000101;
 17'b00001000100100111 : data_comb = 6'b000101;
 17'b00001000100101000 : data_comb = 6'b000100;
 17'b00001000100101001 : data_comb = 6'b111000;
 17'b00001000100101010 : data_comb = 6'b111000;
 17'b00001000100101011 : data_comb = 6'b101000;
 17'b00001000100101100 : data_comb = 6'b000101;
 17'b00001000100101101 : data_comb = 6'b000101;
 17'b00001000100101110 : data_comb = 6'b000101;
 17'b00001000100101111 : data_comb = 6'b000101;
 17'b00001000100110000 : data_comb = 6'b000101;
 17'b00001000100110001 : data_comb = 6'b000101;
 17'b00001000100110010 : data_comb = 6'b000101;
 17'b00001000100110011 : data_comb = 6'b000101;
 17'b00001000100110100 : data_comb = 6'b000101;
 17'b00001000100110101 : data_comb = 6'b000101;
 17'b00001000100110110 : data_comb = 6'b000101;
 17'b00001000100110111 : data_comb = 6'b000101;
 17'b00001000100111000 : data_comb = 6'b000101;
 17'b00001000100111001 : data_comb = 6'b000001;
 17'b00001000100111010 : data_comb = 6'b000001;
 17'b00001000100111011 : data_comb = 6'b000001;
 17'b00001000100111100 : data_comb = 6'b000001;
 17'b00001000100111101 : data_comb = 6'b000001;
 17'b00001000100111110 : data_comb = 6'b000001;
 17'b00001000100111111 : data_comb = 6'b000000;
 17'b00001000101000000 : data_comb = 6'b000000;
 17'b00001000101000001 : data_comb = 6'b000000;
 17'b00001000101000010 : data_comb = 6'b000000;
 17'b00001000101000011 : data_comb = 6'b000000;
 17'b00001000101000100 : data_comb = 6'b000000;
 17'b00001000101000101 : data_comb = 6'b000000;
 17'b00001000101000110 : data_comb = 6'b000000;
 17'b00001000101000111 : data_comb = 6'b010000;
 17'b00001000101001000 : data_comb = 6'b010000;
 17'b00001000101001001 : data_comb = 6'b010000;
 17'b00001000101001010 : data_comb = 6'b010000;
 17'b00001000101001011 : data_comb = 6'b000000;
 17'b00001000101001100 : data_comb = 6'b000000;
 17'b00001000101001101 : data_comb = 6'b000000;
 17'b00001000101001110 : data_comb = 6'b000000;
 17'b00001000101001111 : data_comb = 6'b000000;
 17'b00001000101010000 : data_comb = 6'b010000;
 17'b00001000101010001 : data_comb = 6'b010000;
 17'b00001000101010010 : data_comb = 6'b000000;
 17'b00001000101010011 : data_comb = 6'b000000;
 17'b00001000101010100 : data_comb = 6'b010000;
 17'b00001000101010101 : data_comb = 6'b010000;
 17'b00001000101010110 : data_comb = 6'b010000;
 17'b00001000101010111 : data_comb = 6'b010000;
 17'b00001000101011000 : data_comb = 6'b010000;
 17'b00001000101011001 : data_comb = 6'b010000;
 17'b00001000101011010 : data_comb = 6'b000000;
 17'b00001000101011011 : data_comb = 6'b000000;
 17'b00001000101011100 : data_comb = 6'b010000;
 17'b00001000101011101 : data_comb = 6'b010000;
 17'b00001000101011110 : data_comb = 6'b000000;
 17'b00001000101011111 : data_comb = 6'b000000;
 17'b00001000101100000 : data_comb = 6'b000000;
 17'b00001000101100001 : data_comb = 6'b000000;
 17'b00001000101100010 : data_comb = 6'b000000;
 17'b00001000101100011 : data_comb = 6'b010000;
 17'b00001000101100100 : data_comb = 6'b010000;
 17'b00001000101100101 : data_comb = 6'b010000;
 17'b00001000101100110 : data_comb = 6'b000000;
 17'b00001000101100111 : data_comb = 6'b010000;
 17'b00001000101101000 : data_comb = 6'b010000;
 17'b00001000101101001 : data_comb = 6'b010000;
 17'b00001000101101010 : data_comb = 6'b000000;
 17'b00001000101101011 : data_comb = 6'b000000;
 17'b00001000101101100 : data_comb = 6'b000000;
 17'b00001000101101101 : data_comb = 6'b000000;
 17'b00001000101101110 : data_comb = 6'b000000;
 17'b00001000101101111 : data_comb = 6'b000000;
 17'b00001000101110000 : data_comb = 6'b000000;
 17'b00001000101110001 : data_comb = 6'b000001;
 17'b00001000101110010 : data_comb = 6'b000001;
 17'b00001000101110011 : data_comb = 6'b000001;
 17'b00001000101110100 : data_comb = 6'b000001;
 17'b00001000101110101 : data_comb = 6'b000001;
 17'b00001000101110110 : data_comb = 6'b000001;
 17'b00001000101110111 : data_comb = 6'b000101;
 17'b00001000101111000 : data_comb = 6'b000101;
 17'b00001000101111001 : data_comb = 6'b011000;
 17'b00001000101111010 : data_comb = 6'b010101;
 17'b00001000101111011 : data_comb = 6'b000101;
 17'b00001000101111100 : data_comb = 6'b000101;
 17'b00001000101111101 : data_comb = 6'b000101;
 17'b00001000101111110 : data_comb = 6'b000101;
 17'b00001000101111111 : data_comb = 6'b000101;
 17'b00001000110000000 : data_comb = 6'b000101;
 17'b00001000110000001 : data_comb = 6'b000101;
 17'b00001000110000010 : data_comb = 6'b000101;
 17'b00001000110000011 : data_comb = 6'b000101;
 17'b00001000110000100 : data_comb = 6'b000101;
 17'b00001000110000101 : data_comb = 6'b000101;
 17'b00001000110000110 : data_comb = 6'b000101;
 17'b00001000110000111 : data_comb = 6'b000101;
 17'b00001000110001000 : data_comb = 6'b000001;
 17'b00001000110001001 : data_comb = 6'b000001;
 17'b00001000110001010 : data_comb = 6'b000001;
 17'b00001000110001011 : data_comb = 6'b000001;
 17'b00001000110001100 : data_comb = 6'b000001;
 17'b00001000110001101 : data_comb = 6'b000001;
 17'b00001000110001110 : data_comb = 6'b000001;
 17'b00001000110001111 : data_comb = 6'b000001;
 17'b00001000110010000 : data_comb = 6'b000001;
 17'b00001000110010001 : data_comb = 6'b000001;
 17'b00001000110010010 : data_comb = 6'b000000;
 17'b00001000110010011 : data_comb = 6'b000000;
 17'b00001000110010100 : data_comb = 6'b000000;
 17'b00001000110010101 : data_comb = 6'b000000;
 17'b00001000110010110 : data_comb = 6'b000000;
 17'b00001000110010111 : data_comb = 6'b000000;
 17'b00001000110011000 : data_comb = 6'b000000;
 17'b00001000110011001 : data_comb = 6'b010000;
 17'b00001000110011010 : data_comb = 6'b010000;
 17'b00001000110011011 : data_comb = 6'b000000;
 17'b00001000110011100 : data_comb = 6'b000000;
 17'b00001000110011101 : data_comb = 6'b000000;
 17'b00001000110011110 : data_comb = 6'b000000;
 17'b00001000110011111 : data_comb = 6'b010000;
 17'b00001000110100000 : data_comb = 6'b010000;
 17'b00001000110100001 : data_comb = 6'b010000;
 17'b00001000110100010 : data_comb = 6'b010000;
 17'b00001000110100011 : data_comb = 6'b000000;
 17'b00001000110100100 : data_comb = 6'b000000;
 17'b00001000110100101 : data_comb = 6'b000000;
 17'b00001000110100110 : data_comb = 6'b000000;
 17'b00001000110100111 : data_comb = 6'b000000;
 17'b00001000110101000 : data_comb = 6'b000000;
 17'b00001000110101001 : data_comb = 6'b000000;
 17'b00001000110101010 : data_comb = 6'b000000;
 17'b00001000110101011 : data_comb = 6'b000000;
 17'b00001000110101100 : data_comb = 6'b000000;
 17'b00001000110101101 : data_comb = 6'b000000;
 17'b00001000110101110 : data_comb = 6'b000000;
 17'b00001000110101111 : data_comb = 6'b000000;
 17'b00001000110110000 : data_comb = 6'b000000;
 17'b00001000110110001 : data_comb = 6'b000000;
 17'b00001000110110010 : data_comb = 6'b000000;
 17'b00001000110110011 : data_comb = 6'b000000;
 17'b00001000110110100 : data_comb = 6'b000000;
 17'b00001000110110101 : data_comb = 6'b000000;
 17'b00001000110110110 : data_comb = 6'b000000;
 17'b00001000110110111 : data_comb = 6'b000000;
 17'b00001000110111000 : data_comb = 6'b000000;
 17'b00001000110111001 : data_comb = 6'b000000;
 17'b00001000110111010 : data_comb = 6'b000000;
 17'b00001000110111011 : data_comb = 6'b000000;
 17'b00001000110111100 : data_comb = 6'b000000;
 17'b00001000110111101 : data_comb = 6'b000000;
 17'b00001000110111110 : data_comb = 6'b000000;
 17'b00001000110111111 : data_comb = 6'b000000;
 17'b00001000111000000 : data_comb = 6'b000001;
 17'b00001000111000001 : data_comb = 6'b000001;
 17'b00001000111000010 : data_comb = 6'b000001;
 17'b00001000111000011 : data_comb = 6'b000001;
 17'b00001000111000100 : data_comb = 6'b000001;
 17'b00001000111000101 : data_comb = 6'b000001;
 17'b00001000111000110 : data_comb = 6'b000001;
 17'b00001000111000111 : data_comb = 6'b000001;
 17'b00001000111001000 : data_comb = 6'b000101;
 17'b00001000111001001 : data_comb = 6'b000101;
 17'b00001000111001010 : data_comb = 6'b000101;
 17'b00001000111001011 : data_comb = 6'b000101;
 17'b00001000111001100 : data_comb = 6'b000101;
 17'b00001000111001101 : data_comb = 6'b000101;
 17'b00001000111001110 : data_comb = 6'b000101;
 17'b00001000111001111 : data_comb = 6'b000101;
 17'b00001000111010000 : data_comb = 6'b000101;
 17'b00001000111010001 : data_comb = 6'b000101;
 17'b00001000111010010 : data_comb = 6'b000101;
 17'b00001000111010011 : data_comb = 6'b000101;
 17'b00001000111010100 : data_comb = 6'b000101;
 17'b00001000111010101 : data_comb = 6'b000101;
 17'b00001000111010110 : data_comb = 6'b000101;
 17'b00001000111010111 : data_comb = 6'b000101;
 17'b00001000111011000 : data_comb = 6'b000001;
 17'b00001000111011001 : data_comb = 6'b000001;
 17'b00001000111011010 : data_comb = 6'b000001;
 17'b00001000111011011 : data_comb = 6'b000001;
 17'b00001000111011100 : data_comb = 6'b000001;
 17'b00001000111011101 : data_comb = 6'b000001;
 17'b00001000111011110 : data_comb = 6'b000001;
 17'b00001000111011111 : data_comb = 6'b000001;
 17'b00001000111100000 : data_comb = 6'b000001;
 17'b00001000111100001 : data_comb = 6'b000001;
 17'b00001000111100010 : data_comb = 6'b000000;
 17'b00001000111100011 : data_comb = 6'b000000;
 17'b00001000111100100 : data_comb = 6'b000000;
 17'b00001000111100101 : data_comb = 6'b000000;
 17'b00001000111100110 : data_comb = 6'b000000;
 17'b00001000111100111 : data_comb = 6'b000000;
 17'b00001000111101000 : data_comb = 6'b000000;
 17'b00001000111101001 : data_comb = 6'b000000;
 17'b00001000111101010 : data_comb = 6'b000000;
 17'b00001000111101011 : data_comb = 6'b000000;
 17'b00001000111101100 : data_comb = 6'b000000;
 17'b00001000111101101 : data_comb = 6'b000000;
 17'b00001000111101110 : data_comb = 6'b000000;
 17'b00001000111101111 : data_comb = 6'b000000;
 17'b00001000111110000 : data_comb = 6'b000000;
 17'b00001000111110001 : data_comb = 6'b000000;
 17'b00001000111110010 : data_comb = 6'b000000;
 17'b00001000111110011 : data_comb = 6'b000000;
 17'b00001000111110100 : data_comb = 6'b000000;
 17'b00001000111110101 : data_comb = 6'b000000;
 17'b00001000111110110 : data_comb = 6'b000000;
 17'b00001000111110111 : data_comb = 6'b000000;
 17'b00001000111111000 : data_comb = 6'b000000;
 17'b00001000111111001 : data_comb = 6'b000000;
 17'b00001000111111010 : data_comb = 6'b000000;
 17'b00001000111111011 : data_comb = 6'b000000;
 17'b00001000111111100 : data_comb = 6'b000000;
 17'b00001000111111101 : data_comb = 6'b000000;
 17'b00001000111111110 : data_comb = 6'b000000;
 17'b00001000111111111 : data_comb = 6'b000000;
 17'b00001001000000000 : data_comb = 6'b000000;
 17'b00001001000000001 : data_comb = 6'b000000;
 17'b00001001000000010 : data_comb = 6'b000000;
 17'b00001001000000011 : data_comb = 6'b000000;
 17'b00001001000000100 : data_comb = 6'b000000;
 17'b00001001000000101 : data_comb = 6'b000000;
 17'b00001001000000110 : data_comb = 6'b000000;
 17'b00001001000000111 : data_comb = 6'b000000;
 17'b00001001000001000 : data_comb = 6'b000000;
 17'b00001001000001001 : data_comb = 6'b000000;
 17'b00001001000001010 : data_comb = 6'b000000;
 17'b00001001000001011 : data_comb = 6'b000000;
 17'b00001001000001100 : data_comb = 6'b000000;
 17'b00001001000001101 : data_comb = 6'b000000;
 17'b00001001000001110 : data_comb = 6'b000001;
 17'b00001001000001111 : data_comb = 6'b000001;
 17'b00001001000010000 : data_comb = 6'b000001;
 17'b00001001000010001 : data_comb = 6'b000001;
 17'b00001001000010010 : data_comb = 6'b000001;
 17'b00001001000010011 : data_comb = 6'b000001;
 17'b00001001000010100 : data_comb = 6'b000001;
 17'b00001001000010101 : data_comb = 6'b000001;
 17'b00001001000010110 : data_comb = 6'b000001;
 17'b00001001000010111 : data_comb = 6'b000001;
 17'b00001001000011000 : data_comb = 6'b000001;
 17'b00001001000011001 : data_comb = 6'b000101;
 17'b00001001000011010 : data_comb = 6'b000101;
 17'b00001001000011011 : data_comb = 6'b000101;
 17'b00001001000011100 : data_comb = 6'b000101;
 17'b00001001000011101 : data_comb = 6'b000101;
 17'b00001001000011110 : data_comb = 6'b000101;
 17'b00001001000011111 : data_comb = 6'b000101;
 17'b00001001000100000 : data_comb = 6'b000101;
 17'b00001001000100001 : data_comb = 6'b000101;
 17'b00001001000100010 : data_comb = 6'b000101;
 17'b00001001000100011 : data_comb = 6'b000101;
 17'b00001001000100100 : data_comb = 6'b000101;
 17'b00001001000100101 : data_comb = 6'b000101;
 17'b00001001000100110 : data_comb = 6'b000101;
 17'b00001001000100111 : data_comb = 6'b000101;
 17'b00001001000101000 : data_comb = 6'b000001;
 17'b00001001000101001 : data_comb = 6'b000001;
 17'b00001001000101010 : data_comb = 6'b000001;
 17'b00001001000101011 : data_comb = 6'b000001;
 17'b00001001000101100 : data_comb = 6'b000001;
 17'b00001001000101101 : data_comb = 6'b000001;
 17'b00001001000101110 : data_comb = 6'b000001;
 17'b00001001000101111 : data_comb = 6'b000001;
 17'b00001001000110000 : data_comb = 6'b000001;
 17'b00001001000110001 : data_comb = 6'b000001;
 17'b00001001000110010 : data_comb = 6'b000001;
 17'b00001001000110011 : data_comb = 6'b000001;
 17'b00001001000110100 : data_comb = 6'b000001;
 17'b00001001000110101 : data_comb = 6'b000001;
 17'b00001001000110110 : data_comb = 6'b000001;
 17'b00001001000110111 : data_comb = 6'b000000;
 17'b00001001000111000 : data_comb = 6'b000000;
 17'b00001001000111001 : data_comb = 6'b000000;
 17'b00001001000111010 : data_comb = 6'b000000;
 17'b00001001000111011 : data_comb = 6'b000000;
 17'b00001001000111100 : data_comb = 6'b000000;
 17'b00001001000111101 : data_comb = 6'b000000;
 17'b00001001000111110 : data_comb = 6'b000000;
 17'b00001001000111111 : data_comb = 6'b000000;
 17'b00001001001000000 : data_comb = 6'b000000;
 17'b00001001001000001 : data_comb = 6'b000000;
 17'b00001001001000010 : data_comb = 6'b000000;
 17'b00001001001000011 : data_comb = 6'b000000;
 17'b00001001001000100 : data_comb = 6'b000000;
 17'b00001001001000101 : data_comb = 6'b000000;
 17'b00001001001000110 : data_comb = 6'b000000;
 17'b00001001001000111 : data_comb = 6'b000000;
 17'b00001001001001000 : data_comb = 6'b000000;
 17'b00001001001001001 : data_comb = 6'b000000;
 17'b00001001001001010 : data_comb = 6'b000000;
 17'b00001001001001011 : data_comb = 6'b000000;
 17'b00001001001001100 : data_comb = 6'b000000;
 17'b00001001001001101 : data_comb = 6'b000000;
 17'b00001001001001110 : data_comb = 6'b000000;
 17'b00001001001001111 : data_comb = 6'b000000;
 17'b00001001001010000 : data_comb = 6'b000000;
 17'b00001001001010001 : data_comb = 6'b000000;
 17'b00001001001010010 : data_comb = 6'b000000;
 17'b00001001001010011 : data_comb = 6'b000000;
 17'b00001001001010100 : data_comb = 6'b000000;
 17'b00001001001010101 : data_comb = 6'b000000;
 17'b00001001001010110 : data_comb = 6'b000000;
 17'b00001001001010111 : data_comb = 6'b000000;
 17'b00001001001011000 : data_comb = 6'b000000;
 17'b00001001001011001 : data_comb = 6'b000000;
 17'b00001001001011010 : data_comb = 6'b000000;
 17'b00001001001011011 : data_comb = 6'b000001;
 17'b00001001001011100 : data_comb = 6'b000001;
 17'b00001001001011101 : data_comb = 6'b000001;
 17'b00001001001011110 : data_comb = 6'b000001;
 17'b00001001001011111 : data_comb = 6'b000001;
 17'b00001001001100000 : data_comb = 6'b000001;
 17'b00001001001100001 : data_comb = 6'b000001;
 17'b00001001001100010 : data_comb = 6'b000001;
 17'b00001001001100011 : data_comb = 6'b000001;
 17'b00001001001100100 : data_comb = 6'b000001;
 17'b00001001001100101 : data_comb = 6'b000001;
 17'b00001001001100110 : data_comb = 6'b000001;
 17'b00001001001100111 : data_comb = 6'b000001;
 17'b00001001001101000 : data_comb = 6'b000101;
 17'b00001001001101001 : data_comb = 6'b000101;
 17'b00001001001101010 : data_comb = 6'b000101;
 17'b00001001001101011 : data_comb = 6'b000101;
 17'b00001001001101100 : data_comb = 6'b000101;
 17'b00001001001101101 : data_comb = 6'b000101;
 17'b00001001001101110 : data_comb = 6'b000101;
 17'b00001001001101111 : data_comb = 6'b000101;
 17'b00001001001110000 : data_comb = 6'b000101;
 17'b00001001001110001 : data_comb = 6'b000101;
 17'b00001001001110010 : data_comb = 6'b000101;
 17'b00001001001110011 : data_comb = 6'b000101;
 17'b00001001001110100 : data_comb = 6'b000101;
 17'b00001001001110101 : data_comb = 6'b000101;
 17'b00001001001110110 : data_comb = 6'b000101;
 17'b00001001001110111 : data_comb = 6'b000101;
 17'b00001001001111000 : data_comb = 6'b000001;
 17'b00001001001111001 : data_comb = 6'b000001;
 17'b00001001001111010 : data_comb = 6'b000001;
 17'b00001001001111011 : data_comb = 6'b000001;
 17'b00001001001111100 : data_comb = 6'b000001;
 17'b00001001001111101 : data_comb = 6'b000001;
 17'b00001001001111110 : data_comb = 6'b000001;
 17'b00001001001111111 : data_comb = 6'b000001;
 17'b00001001010000000 : data_comb = 6'b000001;
 17'b00001001010000001 : data_comb = 6'b000001;
 17'b00001001010000010 : data_comb = 6'b000001;
 17'b00001001010000011 : data_comb = 6'b000001;
 17'b00001001010000100 : data_comb = 6'b000001;
 17'b00001001010000101 : data_comb = 6'b000001;
 17'b00001001010000110 : data_comb = 6'b000001;
 17'b00001001010000111 : data_comb = 6'b000001;
 17'b00001001010001000 : data_comb = 6'b000001;
 17'b00001001010001001 : data_comb = 6'b000001;
 17'b00001001010001010 : data_comb = 6'b000001;
 17'b00001001010001011 : data_comb = 6'b000001;
 17'b00001001010001100 : data_comb = 6'b000001;
 17'b00001001010001101 : data_comb = 6'b000001;
 17'b00001001010001110 : data_comb = 6'b000001;
 17'b00001001010001111 : data_comb = 6'b000001;
 17'b00001001010010000 : data_comb = 6'b000001;
 17'b00001001010010001 : data_comb = 6'b000001;
 17'b00001001010010010 : data_comb = 6'b000001;
 17'b00001001010010011 : data_comb = 6'b000001;
 17'b00001001010010100 : data_comb = 6'b000001;
 17'b00001001010010101 : data_comb = 6'b000001;
 17'b00001001010010110 : data_comb = 6'b000001;
 17'b00001001010010111 : data_comb = 6'b000001;
 17'b00001001010011000 : data_comb = 6'b000001;
 17'b00001001010011001 : data_comb = 6'b000001;
 17'b00001001010011010 : data_comb = 6'b000001;
 17'b00001001010011011 : data_comb = 6'b000001;
 17'b00001001010011100 : data_comb = 6'b000001;
 17'b00001001010011101 : data_comb = 6'b000001;
 17'b00001001010011110 : data_comb = 6'b000001;
 17'b00001001010011111 : data_comb = 6'b000001;
 17'b00001001010100000 : data_comb = 6'b000001;
 17'b00001001010100001 : data_comb = 6'b000001;
 17'b00001001010100010 : data_comb = 6'b000001;
 17'b00001001010100011 : data_comb = 6'b000001;
 17'b00001001010100100 : data_comb = 6'b000001;
 17'b00001001010100101 : data_comb = 6'b000001;
 17'b00001001010100110 : data_comb = 6'b000001;
 17'b00001001010100111 : data_comb = 6'b000001;
 17'b00001001010101000 : data_comb = 6'b000001;
 17'b00001001010101001 : data_comb = 6'b000001;
 17'b00001001010101010 : data_comb = 6'b000001;
 17'b00001001010101011 : data_comb = 6'b000001;
 17'b00001001010101100 : data_comb = 6'b000001;
 17'b00001001010101101 : data_comb = 6'b000001;
 17'b00001001010101110 : data_comb = 6'b000001;
 17'b00001001010101111 : data_comb = 6'b000001;
 17'b00001001010110000 : data_comb = 6'b000001;
 17'b00001001010110001 : data_comb = 6'b000001;
 17'b00001001010110010 : data_comb = 6'b000001;
 17'b00001001010110011 : data_comb = 6'b000001;
 17'b00001001010110100 : data_comb = 6'b000001;
 17'b00001001010110101 : data_comb = 6'b000001;
 17'b00001001010110110 : data_comb = 6'b000001;
 17'b00001001010110111 : data_comb = 6'b000001;
 17'b00001001010111000 : data_comb = 6'b000101;
 17'b00001001010111001 : data_comb = 6'b000101;
 17'b00001001010111010 : data_comb = 6'b000101;
 17'b00001001010111011 : data_comb = 6'b000101;
 17'b00001001010111100 : data_comb = 6'b000101;
 17'b00001001010111101 : data_comb = 6'b000101;
 17'b00001001010111110 : data_comb = 6'b000101;
 17'b00001001010111111 : data_comb = 6'b000101;
    default: data_comb = 6'b0;
    endcase
end
endmodule